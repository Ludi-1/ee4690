module toplevel #(
    parameter MATRIX_DIM = 64,
    parameter INPUT_WIDTH = 8,
    parameter OUTPUT_WIDTH = 20,
)

(
    input CLK,
    input rst
);

always @ (posedge CLK) begin
    
end



endmodule