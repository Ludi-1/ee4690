module fc (
    input CLK,
    
)

endmodule