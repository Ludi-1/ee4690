module conv_layer #(
    parameter input_channels = 1, // DO NOT CHANGE for now, others are unsupported.
    parameter input_size = 28, // Size of the input image. Size is symmetric.
    parameter output_channels = 16 // Amount of output channels.
) (
    input clk, reset, i_write_enable, i_data
);

endmodule