module layer_3_conv #(
    parameter INPUT_DIM = 28,   //28x28
    parameter OUTPUT_DIM = 10,
    parameter KERNEL_DIM = 3,
    parameter INPUT_CHANNELS = 1,
    parameter OUTPUT_CHANNELS = 2,
    parameter DATATYPE_SIZE = 1
) (
    input clk,
    input reset,

    input i_we,
    input [DATATYPE_SIZE-1:0] i_data [INPUT_CHANNELS-1:0],

    output [DATATYPE_SIZE-1:0] o_data [OUTPUT_CHANNELS-1:0],
    output o_we
);

localparam TEMP_SIZE = INPUT_CHANNELS * OUTPUT_CHANNELS * (KERNAL_DIM ** 2);

reg window [INPUT_CHANNELS-1:0][KERNAL_DIM**2-1:0];
reg temp [TEMP_SIZE-1:0];

ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[0]),
                        .o_data(window[0]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[1]),
                        .o_data(window[1]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[2]),
                        .o_data(window[2]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[3]),
                        .o_data(window[3]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[4]),
                        .o_data(window[4]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[5]),
                        .o_data(window[5]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[6]),
                        .o_data(window[6]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[7]),
                        .o_data(window[7]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[8]),
                        .o_data(window[8]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[9]),
                        .o_data(window[9]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[10]),
                        .o_data(window[10]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[11]),
                        .o_data(window[11]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[12]),
                        .o_data(window[12]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[13]),
                        .o_data(window[13]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[14]),
                        .o_data(window[14]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[15]),
                        .o_data(window[15]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[16]),
                        .o_data(window[16]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[17]),
                        .o_data(window[17]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[18]),
                        .o_data(window[18]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[19]),
                        .o_data(window[19]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[20]),
                        .o_data(window[20]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[21]),
                        .o_data(window[21]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[22]),
                        .o_data(window[22]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[23]),
                        .o_data(window[23]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[24]),
                        .o_data(window[24]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[25]),
                        .o_data(window[25]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[26]),
                        .o_data(window[26]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[27]),
                        .o_data(window[27]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[28]),
                        .o_data(window[28]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[29]),
                        .o_data(window[29]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[30]),
                        .o_data(window[30]),
                    );
ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[31]),
                        .o_data(window[31]),
                    );

# ibuf_conv #(
#     .img_width(INPUT_DIM),
#     .kernel_dim(KERNEL_DIM),
# ) ibuf (
#     .clk(clk),
#     .i_we(i_we),
#     .i_data(i_data[%INPUT_C%]),
#     .o_data(window[%INPUT_C%]),
# );

assign temp[0] = window[0][0];
assign temp[1] = ~window[0][1];
assign temp[2] = window[0][2];
assign temp[3] = window[0][3];
assign temp[4] = ~window[0][4];
assign temp[5] = window[0][5];
assign temp[6] = ~window[0][6];
assign temp[7] = ~window[0][7];
assign temp[8] = window[0][8];
assign temp[32] = ~window[1][0];
assign temp[33] = ~window[1][1];
assign temp[34] = ~window[1][2];
assign temp[35] = window[1][3];
assign temp[36] = ~window[1][4];
assign temp[37] = window[1][5];
assign temp[38] = window[1][6];
assign temp[39] = ~window[1][7];
assign temp[40] = ~window[1][8];
assign temp[64] = ~window[2][0];
assign temp[65] = ~window[2][1];
assign temp[66] = ~window[2][2];
assign temp[67] = window[2][3];
assign temp[68] = ~window[2][4];
assign temp[69] = ~window[2][5];
assign temp[70] = window[2][6];
assign temp[71] = ~window[2][7];
assign temp[72] = ~window[2][8];
assign temp[96] = window[3][0];
assign temp[97] = ~window[3][1];
assign temp[98] = window[3][2];
assign temp[99] = window[3][3];
assign temp[100] = ~window[3][4];
assign temp[101] = window[3][5];
assign temp[102] = window[3][6];
assign temp[103] = ~window[3][7];
assign temp[104] = window[3][8];
assign temp[128] = window[4][0];
assign temp[129] = window[4][1];
assign temp[130] = ~window[4][2];
assign temp[131] = ~window[4][3];
assign temp[132] = ~window[4][4];
assign temp[133] = ~window[4][5];
assign temp[134] = ~window[4][6];
assign temp[135] = ~window[4][7];
assign temp[136] = ~window[4][8];
assign temp[160] = window[5][0];
assign temp[161] = ~window[5][1];
assign temp[162] = window[5][2];
assign temp[163] = window[5][3];
assign temp[164] = ~window[5][4];
assign temp[165] = window[5][5];
assign temp[166] = ~window[5][6];
assign temp[167] = ~window[5][7];
assign temp[168] = window[5][8];
assign temp[192] = window[6][0];
assign temp[193] = window[6][1];
assign temp[194] = ~window[6][2];
assign temp[195] = ~window[6][3];
assign temp[196] = window[6][4];
assign temp[197] = ~window[6][5];
assign temp[198] = window[6][6];
assign temp[199] = ~window[6][7];
assign temp[200] = ~window[6][8];
assign temp[224] = window[7][0];
assign temp[225] = ~window[7][1];
assign temp[226] = window[7][2];
assign temp[227] = window[7][3];
assign temp[228] = ~window[7][4];
assign temp[229] = window[7][5];
assign temp[230] = ~window[7][6];
assign temp[231] = ~window[7][7];
assign temp[232] = window[7][8];
assign temp[256] = ~window[8][0];
assign temp[257] = ~window[8][1];
assign temp[258] = window[8][2];
assign temp[259] = ~window[8][3];
assign temp[260] = window[8][4];
assign temp[261] = window[8][5];
assign temp[262] = ~window[8][6];
assign temp[263] = window[8][7];
assign temp[264] = ~window[8][8];
assign temp[288] = ~window[9][0];
assign temp[289] = ~window[9][1];
assign temp[290] = window[9][2];
assign temp[291] = window[9][3];
assign temp[292] = ~window[9][4];
assign temp[293] = ~window[9][5];
assign temp[294] = window[9][6];
assign temp[295] = window[9][7];
assign temp[296] = window[9][8];
assign temp[320] = window[10][0];
assign temp[321] = ~window[10][1];
assign temp[322] = ~window[10][2];
assign temp[323] = window[10][3];
assign temp[324] = ~window[10][4];
assign temp[325] = ~window[10][5];
assign temp[326] = ~window[10][6];
assign temp[327] = ~window[10][7];
assign temp[328] = ~window[10][8];
assign temp[352] = window[11][0];
assign temp[353] = ~window[11][1];
assign temp[354] = ~window[11][2];
assign temp[355] = window[11][3];
assign temp[356] = ~window[11][4];
assign temp[357] = ~window[11][5];
assign temp[358] = ~window[11][6];
assign temp[359] = ~window[11][7];
assign temp[360] = ~window[11][8];
assign temp[384] = ~window[12][0];
assign temp[385] = window[12][1];
assign temp[386] = ~window[12][2];
assign temp[387] = window[12][3];
assign temp[388] = window[12][4];
assign temp[389] = window[12][5];
assign temp[390] = window[12][6];
assign temp[391] = window[12][7];
assign temp[392] = ~window[12][8];
assign temp[416] = window[13][0];
assign temp[417] = window[13][1];
assign temp[418] = ~window[13][2];
assign temp[419] = window[13][3];
assign temp[420] = window[13][4];
assign temp[421] = ~window[13][5];
assign temp[422] = window[13][6];
assign temp[423] = ~window[13][7];
assign temp[424] = ~window[13][8];
assign temp[448] = ~window[14][0];
assign temp[449] = ~window[14][1];
assign temp[450] = ~window[14][2];
assign temp[451] = window[14][3];
assign temp[452] = ~window[14][4];
assign temp[453] = window[14][5];
assign temp[454] = ~window[14][6];
assign temp[455] = window[14][7];
assign temp[456] = window[14][8];
assign temp[480] = window[15][0];
assign temp[481] = window[15][1];
assign temp[482] = ~window[15][2];
assign temp[483] = ~window[15][3];
assign temp[484] = window[15][4];
assign temp[485] = ~window[15][5];
assign temp[486] = window[15][6];
assign temp[487] = ~window[15][7];
assign temp[488] = ~window[15][8];
assign temp[512] = window[16][0];
assign temp[513] = window[16][1];
assign temp[514] = window[16][2];
assign temp[515] = ~window[16][3];
assign temp[516] = window[16][4];
assign temp[517] = window[16][5];
assign temp[518] = ~window[16][6];
assign temp[519] = window[16][7];
assign temp[520] = window[16][8];
assign temp[544] = ~window[17][0];
assign temp[545] = ~window[17][1];
assign temp[546] = ~window[17][2];
assign temp[547] = window[17][3];
assign temp[548] = ~window[17][4];
assign temp[549] = window[17][5];
assign temp[550] = window[17][6];
assign temp[551] = window[17][7];
assign temp[552] = window[17][8];
assign temp[576] = ~window[18][0];
assign temp[577] = window[18][1];
assign temp[578] = ~window[18][2];
assign temp[579] = ~window[18][3];
assign temp[580] = window[18][4];
assign temp[581] = ~window[18][5];
assign temp[582] = window[18][6];
assign temp[583] = window[18][7];
assign temp[584] = ~window[18][8];
assign temp[608] = window[19][0];
assign temp[609] = ~window[19][1];
assign temp[610] = ~window[19][2];
assign temp[611] = ~window[19][3];
assign temp[612] = ~window[19][4];
assign temp[613] = ~window[19][5];
assign temp[614] = window[19][6];
assign temp[615] = ~window[19][7];
assign temp[616] = window[19][8];
assign temp[640] = ~window[20][0];
assign temp[641] = ~window[20][1];
assign temp[642] = ~window[20][2];
assign temp[643] = window[20][3];
assign temp[644] = ~window[20][4];
assign temp[645] = window[20][5];
assign temp[646] = ~window[20][6];
assign temp[647] = ~window[20][7];
assign temp[648] = window[20][8];
assign temp[672] = window[21][0];
assign temp[673] = ~window[21][1];
assign temp[674] = ~window[21][2];
assign temp[675] = window[21][3];
assign temp[676] = ~window[21][4];
assign temp[677] = ~window[21][5];
assign temp[678] = ~window[21][6];
assign temp[679] = ~window[21][7];
assign temp[680] = window[21][8];
assign temp[704] = window[22][0];
assign temp[705] = window[22][1];
assign temp[706] = window[22][2];
assign temp[707] = ~window[22][3];
assign temp[708] = window[22][4];
assign temp[709] = ~window[22][5];
assign temp[710] = ~window[22][6];
assign temp[711] = window[22][7];
assign temp[712] = ~window[22][8];
assign temp[736] = ~window[23][0];
assign temp[737] = ~window[23][1];
assign temp[738] = window[23][2];
assign temp[739] = window[23][3];
assign temp[740] = ~window[23][4];
assign temp[741] = window[23][5];
assign temp[742] = window[23][6];
assign temp[743] = ~window[23][7];
assign temp[744] = window[23][8];
assign temp[768] = ~window[24][0];
assign temp[769] = ~window[24][1];
assign temp[770] = ~window[24][2];
assign temp[771] = window[24][3];
assign temp[772] = ~window[24][4];
assign temp[773] = window[24][5];
assign temp[774] = window[24][6];
assign temp[775] = ~window[24][7];
assign temp[776] = ~window[24][8];
assign temp[800] = ~window[25][0];
assign temp[801] = ~window[25][1];
assign temp[802] = window[25][2];
assign temp[803] = window[25][3];
assign temp[804] = window[25][4];
assign temp[805] = window[25][5];
assign temp[806] = window[25][6];
assign temp[807] = window[25][7];
assign temp[808] = window[25][8];
assign temp[832] = window[26][0];
assign temp[833] = ~window[26][1];
assign temp[834] = ~window[26][2];
assign temp[835] = window[26][3];
assign temp[836] = ~window[26][4];
assign temp[837] = ~window[26][5];
assign temp[838] = window[26][6];
assign temp[839] = ~window[26][7];
assign temp[840] = window[26][8];
assign temp[864] = window[27][0];
assign temp[865] = ~window[27][1];
assign temp[866] = window[27][2];
assign temp[867] = window[27][3];
assign temp[868] = window[27][4];
assign temp[869] = window[27][5];
assign temp[870] = ~window[27][6];
assign temp[871] = ~window[27][7];
assign temp[872] = window[27][8];
assign temp[896] = ~window[28][0];
assign temp[897] = window[28][1];
assign temp[898] = window[28][2];
assign temp[899] = ~window[28][3];
assign temp[900] = window[28][4];
assign temp[901] = ~window[28][5];
assign temp[902] = window[28][6];
assign temp[903] = window[28][7];
assign temp[904] = ~window[28][8];
assign temp[928] = window[29][0];
assign temp[929] = ~window[29][1];
assign temp[930] = ~window[29][2];
assign temp[931] = window[29][3];
assign temp[932] = ~window[29][4];
assign temp[933] = ~window[29][5];
assign temp[934] = ~window[29][6];
assign temp[935] = ~window[29][7];
assign temp[936] = ~window[29][8];
assign temp[960] = ~window[30][0];
assign temp[961] = window[30][1];
assign temp[962] = window[30][2];
assign temp[963] = ~window[30][3];
assign temp[964] = window[30][4];
assign temp[965] = window[30][5];
assign temp[966] = window[30][6];
assign temp[967] = window[30][7];
assign temp[968] = window[30][8];
assign temp[992] = ~window[31][0];
assign temp[993] = ~window[31][1];
assign temp[994] = ~window[31][2];
assign temp[995] = window[31][3];
assign temp[996] = window[31][4];
assign temp[997] = ~window[31][5];
assign temp[998] = window[31][6];
assign temp[999] = ~window[31][7];
assign temp[1000] = ~window[31][8];
assign temp[32] = ~window[0][0];
assign temp[33] = window[0][1];
assign temp[34] = ~window[0][2];
assign temp[35] = ~window[0][3];
assign temp[36] = ~window[0][4];
assign temp[37] = window[0][5];
assign temp[38] = ~window[0][6];
assign temp[39] = ~window[0][7];
assign temp[40] = window[0][8];
assign temp[64] = window[1][0];
assign temp[65] = ~window[1][1];
assign temp[66] = ~window[1][2];
assign temp[67] = ~window[1][3];
assign temp[68] = ~window[1][4];
assign temp[69] = window[1][5];
assign temp[70] = window[1][6];
assign temp[71] = window[1][7];
assign temp[72] = window[1][8];
assign temp[96] = ~window[2][0];
assign temp[97] = window[2][1];
assign temp[98] = ~window[2][2];
assign temp[99] = window[2][3];
assign temp[100] = window[2][4];
assign temp[101] = window[2][5];
assign temp[102] = window[2][6];
assign temp[103] = window[2][7];
assign temp[104] = window[2][8];
assign temp[128] = window[3][0];
assign temp[129] = ~window[3][1];
assign temp[130] = ~window[3][2];
assign temp[131] = window[3][3];
assign temp[132] = window[3][4];
assign temp[133] = window[3][5];
assign temp[134] = window[3][6];
assign temp[135] = window[3][7];
assign temp[136] = window[3][8];
assign temp[160] = ~window[4][0];
assign temp[161] = ~window[4][1];
assign temp[162] = window[4][2];
assign temp[163] = window[4][3];
assign temp[164] = window[4][4];
assign temp[165] = window[4][5];
assign temp[166] = window[4][6];
assign temp[167] = ~window[4][7];
assign temp[168] = ~window[4][8];
assign temp[192] = ~window[5][0];
assign temp[193] = ~window[5][1];
assign temp[194] = ~window[5][2];
assign temp[195] = ~window[5][3];
assign temp[196] = window[5][4];
assign temp[197] = ~window[5][5];
assign temp[198] = ~window[5][6];
assign temp[199] = ~window[5][7];
assign temp[200] = ~window[5][8];
assign temp[224] = window[6][0];
assign temp[225] = ~window[6][1];
assign temp[226] = ~window[6][2];
assign temp[227] = window[6][3];
assign temp[228] = window[6][4];
assign temp[229] = window[6][5];
assign temp[230] = ~window[6][6];
assign temp[231] = window[6][7];
assign temp[232] = window[6][8];
assign temp[256] = window[7][0];
assign temp[257] = ~window[7][1];
assign temp[258] = ~window[7][2];
assign temp[259] = window[7][3];
assign temp[260] = window[7][4];
assign temp[261] = window[7][5];
assign temp[262] = ~window[7][6];
assign temp[263] = ~window[7][7];
assign temp[264] = ~window[7][8];
assign temp[288] = window[8][0];
assign temp[289] = ~window[8][1];
assign temp[290] = window[8][2];
assign temp[291] = window[8][3];
assign temp[292] = window[8][4];
assign temp[293] = window[8][5];
assign temp[294] = window[8][6];
assign temp[295] = window[8][7];
assign temp[296] = window[8][8];
assign temp[320] = window[9][0];
assign temp[321] = window[9][1];
assign temp[322] = ~window[9][2];
assign temp[323] = window[9][3];
assign temp[324] = window[9][4];
assign temp[325] = ~window[9][5];
assign temp[326] = window[9][6];
assign temp[327] = window[9][7];
assign temp[328] = window[9][8];
assign temp[352] = window[10][0];
assign temp[353] = ~window[10][1];
assign temp[354] = ~window[10][2];
assign temp[355] = ~window[10][3];
assign temp[356] = window[10][4];
assign temp[357] = window[10][5];
assign temp[358] = window[10][6];
assign temp[359] = window[10][7];
assign temp[360] = ~window[10][8];
assign temp[384] = ~window[11][0];
assign temp[385] = window[11][1];
assign temp[386] = window[11][2];
assign temp[387] = window[11][3];
assign temp[388] = window[11][4];
assign temp[389] = window[11][5];
assign temp[390] = ~window[11][6];
assign temp[391] = ~window[11][7];
assign temp[392] = ~window[11][8];
assign temp[416] = ~window[12][0];
assign temp[417] = window[12][1];
assign temp[418] = ~window[12][2];
assign temp[419] = ~window[12][3];
assign temp[420] = window[12][4];
assign temp[421] = window[12][5];
assign temp[422] = window[12][6];
assign temp[423] = window[12][7];
assign temp[424] = window[12][8];
assign temp[448] = ~window[13][0];
assign temp[449] = ~window[13][1];
assign temp[450] = window[13][2];
assign temp[451] = window[13][3];
assign temp[452] = window[13][4];
assign temp[453] = ~window[13][5];
assign temp[454] = ~window[13][6];
assign temp[455] = window[13][7];
assign temp[456] = window[13][8];
assign temp[480] = window[14][0];
assign temp[481] = ~window[14][1];
assign temp[482] = window[14][2];
assign temp[483] = window[14][3];
assign temp[484] = window[14][4];
assign temp[485] = window[14][5];
assign temp[486] = ~window[14][6];
assign temp[487] = ~window[14][7];
assign temp[488] = ~window[14][8];
assign temp[512] = window[15][0];
assign temp[513] = window[15][1];
assign temp[514] = ~window[15][2];
assign temp[515] = ~window[15][3];
assign temp[516] = ~window[15][4];
assign temp[517] = ~window[15][5];
assign temp[518] = ~window[15][6];
assign temp[519] = window[15][7];
assign temp[520] = window[15][8];
assign temp[544] = window[16][0];
assign temp[545] = window[16][1];
assign temp[546] = window[16][2];
assign temp[547] = window[16][3];
assign temp[548] = window[16][4];
assign temp[549] = window[16][5];
assign temp[550] = ~window[16][6];
assign temp[551] = ~window[16][7];
assign temp[552] = ~window[16][8];
assign temp[576] = window[17][0];
assign temp[577] = ~window[17][1];
assign temp[578] = ~window[17][2];
assign temp[579] = ~window[17][3];
assign temp[580] = window[17][4];
assign temp[581] = ~window[17][5];
assign temp[582] = window[17][6];
assign temp[583] = window[17][7];
assign temp[584] = window[17][8];
assign temp[608] = window[18][0];
assign temp[609] = window[18][1];
assign temp[610] = window[18][2];
assign temp[611] = ~window[18][3];
assign temp[612] = window[18][4];
assign temp[613] = ~window[18][5];
assign temp[614] = window[18][6];
assign temp[615] = window[18][7];
assign temp[616] = window[18][8];
assign temp[640] = ~window[19][0];
assign temp[641] = ~window[19][1];
assign temp[642] = ~window[19][2];
assign temp[643] = ~window[19][3];
assign temp[644] = ~window[19][4];
assign temp[645] = ~window[19][5];
assign temp[646] = window[19][6];
assign temp[647] = ~window[19][7];
assign temp[648] = ~window[19][8];
assign temp[672] = window[20][0];
assign temp[673] = window[20][1];
assign temp[674] = window[20][2];
assign temp[675] = window[20][3];
assign temp[676] = window[20][4];
assign temp[677] = window[20][5];
assign temp[678] = window[20][6];
assign temp[679] = window[20][7];
assign temp[680] = window[20][8];
assign temp[704] = ~window[21][0];
assign temp[705] = ~window[21][1];
assign temp[706] = ~window[21][2];
assign temp[707] = window[21][3];
assign temp[708] = ~window[21][4];
assign temp[709] = ~window[21][5];
assign temp[710] = ~window[21][6];
assign temp[711] = ~window[21][7];
assign temp[712] = ~window[21][8];
assign temp[736] = ~window[22][0];
assign temp[737] = window[22][1];
assign temp[738] = window[22][2];
assign temp[739] = window[22][3];
assign temp[740] = window[22][4];
assign temp[741] = ~window[22][5];
assign temp[742] = ~window[22][6];
assign temp[743] = ~window[22][7];
assign temp[744] = window[22][8];
assign temp[768] = ~window[23][0];
assign temp[769] = ~window[23][1];
assign temp[770] = window[23][2];
assign temp[771] = window[23][3];
assign temp[772] = ~window[23][4];
assign temp[773] = ~window[23][5];
assign temp[774] = window[23][6];
assign temp[775] = ~window[23][7];
assign temp[776] = ~window[23][8];
assign temp[800] = window[24][0];
assign temp[801] = ~window[24][1];
assign temp[802] = window[24][2];
assign temp[803] = ~window[24][3];
assign temp[804] = window[24][4];
assign temp[805] = window[24][5];
assign temp[806] = window[24][6];
assign temp[807] = window[24][7];
assign temp[808] = window[24][8];
assign temp[832] = window[25][0];
assign temp[833] = ~window[25][1];
assign temp[834] = window[25][2];
assign temp[835] = window[25][3];
assign temp[836] = ~window[25][4];
assign temp[837] = window[25][5];
assign temp[838] = window[25][6];
assign temp[839] = ~window[25][7];
assign temp[840] = window[25][8];
assign temp[864] = ~window[26][0];
assign temp[865] = ~window[26][1];
assign temp[866] = ~window[26][2];
assign temp[867] = ~window[26][3];
assign temp[868] = ~window[26][4];
assign temp[869] = ~window[26][5];
assign temp[870] = window[26][6];
assign temp[871] = ~window[26][7];
assign temp[872] = ~window[26][8];
assign temp[896] = ~window[27][0];
assign temp[897] = window[27][1];
assign temp[898] = ~window[27][2];
assign temp[899] = window[27][3];
assign temp[900] = window[27][4];
assign temp[901] = ~window[27][5];
assign temp[902] = ~window[27][6];
assign temp[903] = ~window[27][7];
assign temp[904] = ~window[27][8];
assign temp[928] = window[28][0];
assign temp[929] = window[28][1];
assign temp[930] = window[28][2];
assign temp[931] = window[28][3];
assign temp[932] = window[28][4];
assign temp[933] = window[28][5];
assign temp[934] = window[28][6];
assign temp[935] = ~window[28][7];
assign temp[936] = window[28][8];
assign temp[960] = ~window[29][0];
assign temp[961] = window[29][1];
assign temp[962] = window[29][2];
assign temp[963] = window[29][3];
assign temp[964] = window[29][4];
assign temp[965] = ~window[29][5];
assign temp[966] = window[29][6];
assign temp[967] = ~window[29][7];
assign temp[968] = ~window[29][8];
assign temp[992] = window[30][0];
assign temp[993] = window[30][1];
assign temp[994] = ~window[30][2];
assign temp[995] = window[30][3];
assign temp[996] = ~window[30][4];
assign temp[997] = ~window[30][5];
assign temp[998] = ~window[30][6];
assign temp[999] = ~window[30][7];
assign temp[1000] = ~window[30][8];
assign temp[1024] = ~window[31][0];
assign temp[1025] = window[31][1];
assign temp[1026] = window[31][2];
assign temp[1027] = window[31][3];
assign temp[1028] = window[31][4];
assign temp[1029] = window[31][5];
assign temp[1030] = window[31][6];
assign temp[1031] = window[31][7];
assign temp[1032] = window[31][8];
assign temp[64] = ~window[0][0];
assign temp[65] = ~window[0][1];
assign temp[66] = ~window[0][2];
assign temp[67] = window[0][3];
assign temp[68] = window[0][4];
assign temp[69] = window[0][5];
assign temp[70] = ~window[0][6];
assign temp[71] = window[0][7];
assign temp[72] = window[0][8];
assign temp[96] = window[1][0];
assign temp[97] = ~window[1][1];
assign temp[98] = window[1][2];
assign temp[99] = window[1][3];
assign temp[100] = window[1][4];
assign temp[101] = ~window[1][5];
assign temp[102] = window[1][6];
assign temp[103] = window[1][7];
assign temp[104] = ~window[1][8];
assign temp[128] = ~window[2][0];
assign temp[129] = ~window[2][1];
assign temp[130] = window[2][2];
assign temp[131] = window[2][3];
assign temp[132] = window[2][4];
assign temp[133] = window[2][5];
assign temp[134] = window[2][6];
assign temp[135] = window[2][7];
assign temp[136] = window[2][8];
assign temp[160] = window[3][0];
assign temp[161] = ~window[3][1];
assign temp[162] = ~window[3][2];
assign temp[163] = window[3][3];
assign temp[164] = window[3][4];
assign temp[165] = window[3][5];
assign temp[166] = ~window[3][6];
assign temp[167] = ~window[3][7];
assign temp[168] = window[3][8];
assign temp[192] = window[4][0];
assign temp[193] = window[4][1];
assign temp[194] = window[4][2];
assign temp[195] = ~window[4][3];
assign temp[196] = window[4][4];
assign temp[197] = window[4][5];
assign temp[198] = ~window[4][6];
assign temp[199] = ~window[4][7];
assign temp[200] = window[4][8];
assign temp[224] = ~window[5][0];
assign temp[225] = window[5][1];
assign temp[226] = ~window[5][2];
assign temp[227] = ~window[5][3];
assign temp[228] = window[5][4];
assign temp[229] = window[5][5];
assign temp[230] = ~window[5][6];
assign temp[231] = ~window[5][7];
assign temp[232] = window[5][8];
assign temp[256] = ~window[6][0];
assign temp[257] = ~window[6][1];
assign temp[258] = ~window[6][2];
assign temp[259] = ~window[6][3];
assign temp[260] = window[6][4];
assign temp[261] = window[6][5];
assign temp[262] = window[6][6];
assign temp[263] = window[6][7];
assign temp[264] = window[6][8];
assign temp[288] = window[7][0];
assign temp[289] = window[7][1];
assign temp[290] = window[7][2];
assign temp[291] = ~window[7][3];
assign temp[292] = window[7][4];
assign temp[293] = window[7][5];
assign temp[294] = ~window[7][6];
assign temp[295] = ~window[7][7];
assign temp[296] = window[7][8];
assign temp[320] = window[8][0];
assign temp[321] = window[8][1];
assign temp[322] = window[8][2];
assign temp[323] = window[8][3];
assign temp[324] = window[8][4];
assign temp[325] = window[8][5];
assign temp[326] = ~window[8][6];
assign temp[327] = window[8][7];
assign temp[328] = window[8][8];
assign temp[352] = ~window[9][0];
assign temp[353] = ~window[9][1];
assign temp[354] = ~window[9][2];
assign temp[355] = ~window[9][3];
assign temp[356] = window[9][4];
assign temp[357] = window[9][5];
assign temp[358] = window[9][6];
assign temp[359] = window[9][7];
assign temp[360] = ~window[9][8];
assign temp[384] = window[10][0];
assign temp[385] = window[10][1];
assign temp[386] = ~window[10][2];
assign temp[387] = window[10][3];
assign temp[388] = ~window[10][4];
assign temp[389] = window[10][5];
assign temp[390] = ~window[10][6];
assign temp[391] = ~window[10][7];
assign temp[392] = ~window[10][8];
assign temp[416] = window[11][0];
assign temp[417] = window[11][1];
assign temp[418] = window[11][2];
assign temp[419] = ~window[11][3];
assign temp[420] = ~window[11][4];
assign temp[421] = window[11][5];
assign temp[422] = ~window[11][6];
assign temp[423] = ~window[11][7];
assign temp[424] = ~window[11][8];
assign temp[448] = ~window[12][0];
assign temp[449] = ~window[12][1];
assign temp[450] = ~window[12][2];
assign temp[451] = window[12][3];
assign temp[452] = ~window[12][4];
assign temp[453] = ~window[12][5];
assign temp[454] = ~window[12][6];
assign temp[455] = window[12][7];
assign temp[456] = ~window[12][8];
assign temp[480] = ~window[13][0];
assign temp[481] = window[13][1];
assign temp[482] = ~window[13][2];
assign temp[483] = ~window[13][3];
assign temp[484] = ~window[13][4];
assign temp[485] = ~window[13][5];
assign temp[486] = ~window[13][6];
assign temp[487] = ~window[13][7];
assign temp[488] = ~window[13][8];
assign temp[512] = window[14][0];
assign temp[513] = window[14][1];
assign temp[514] = ~window[14][2];
assign temp[515] = window[14][3];
assign temp[516] = window[14][4];
assign temp[517] = window[14][5];
assign temp[518] = ~window[14][6];
assign temp[519] = ~window[14][7];
assign temp[520] = ~window[14][8];
assign temp[544] = ~window[15][0];
assign temp[545] = window[15][1];
assign temp[546] = window[15][2];
assign temp[547] = ~window[15][3];
assign temp[548] = ~window[15][4];
assign temp[549] = window[15][5];
assign temp[550] = window[15][6];
assign temp[551] = window[15][7];
assign temp[552] = window[15][8];
assign temp[576] = ~window[16][0];
assign temp[577] = ~window[16][1];
assign temp[578] = window[16][2];
assign temp[579] = ~window[16][3];
assign temp[580] = window[16][4];
assign temp[581] = window[16][5];
assign temp[582] = ~window[16][6];
assign temp[583] = ~window[16][7];
assign temp[584] = window[16][8];
assign temp[608] = ~window[17][0];
assign temp[609] = window[17][1];
assign temp[610] = ~window[17][2];
assign temp[611] = window[17][3];
assign temp[612] = window[17][4];
assign temp[613] = window[17][5];
assign temp[614] = ~window[17][6];
assign temp[615] = ~window[17][7];
assign temp[616] = ~window[17][8];
assign temp[640] = window[18][0];
assign temp[641] = window[18][1];
assign temp[642] = window[18][2];
assign temp[643] = ~window[18][3];
assign temp[644] = window[18][4];
assign temp[645] = ~window[18][5];
assign temp[646] = window[18][6];
assign temp[647] = window[18][7];
assign temp[648] = window[18][8];
assign temp[672] = window[19][0];
assign temp[673] = window[19][1];
assign temp[674] = ~window[19][2];
assign temp[675] = window[19][3];
assign temp[676] = ~window[19][4];
assign temp[677] = ~window[19][5];
assign temp[678] = window[19][6];
assign temp[679] = ~window[19][7];
assign temp[680] = ~window[19][8];
assign temp[704] = ~window[20][0];
assign temp[705] = ~window[20][1];
assign temp[706] = ~window[20][2];
assign temp[707] = window[20][3];
assign temp[708] = window[20][4];
assign temp[709] = window[20][5];
assign temp[710] = window[20][6];
assign temp[711] = window[20][7];
assign temp[712] = window[20][8];
assign temp[736] = ~window[21][0];
assign temp[737] = ~window[21][1];
assign temp[738] = ~window[21][2];
assign temp[739] = ~window[21][3];
assign temp[740] = ~window[21][4];
assign temp[741] = ~window[21][5];
assign temp[742] = ~window[21][6];
assign temp[743] = ~window[21][7];
assign temp[744] = ~window[21][8];
assign temp[768] = window[22][0];
assign temp[769] = window[22][1];
assign temp[770] = window[22][2];
assign temp[771] = ~window[22][3];
assign temp[772] = window[22][4];
assign temp[773] = window[22][5];
assign temp[774] = ~window[22][6];
assign temp[775] = ~window[22][7];
assign temp[776] = ~window[22][8];
assign temp[800] = ~window[23][0];
assign temp[801] = ~window[23][1];
assign temp[802] = ~window[23][2];
assign temp[803] = window[23][3];
assign temp[804] = window[23][4];
assign temp[805] = window[23][5];
assign temp[806] = ~window[23][6];
assign temp[807] = ~window[23][7];
assign temp[808] = window[23][8];
assign temp[832] = window[24][0];
assign temp[833] = ~window[24][1];
assign temp[834] = window[24][2];
assign temp[835] = window[24][3];
assign temp[836] = window[24][4];
assign temp[837] = window[24][5];
assign temp[838] = window[24][6];
assign temp[839] = window[24][7];
assign temp[840] = window[24][8];
assign temp[864] = ~window[25][0];
assign temp[865] = window[25][1];
assign temp[866] = ~window[25][2];
assign temp[867] = window[25][3];
assign temp[868] = window[25][4];
assign temp[869] = window[25][5];
assign temp[870] = ~window[25][6];
assign temp[871] = ~window[25][7];
assign temp[872] = window[25][8];
assign temp[896] = ~window[26][0];
assign temp[897] = ~window[26][1];
assign temp[898] = ~window[26][2];
assign temp[899] = ~window[26][3];
assign temp[900] = window[26][4];
assign temp[901] = window[26][5];
assign temp[902] = window[26][6];
assign temp[903] = ~window[26][7];
assign temp[904] = ~window[26][8];
assign temp[928] = ~window[27][0];
assign temp[929] = window[27][1];
assign temp[930] = window[27][2];
assign temp[931] = ~window[27][3];
assign temp[932] = window[27][4];
assign temp[933] = window[27][5];
assign temp[934] = ~window[27][6];
assign temp[935] = ~window[27][7];
assign temp[936] = ~window[27][8];
assign temp[960] = window[28][0];
assign temp[961] = window[28][1];
assign temp[962] = window[28][2];
assign temp[963] = window[28][3];
assign temp[964] = ~window[28][4];
assign temp[965] = window[28][5];
assign temp[966] = ~window[28][6];
assign temp[967] = ~window[28][7];
assign temp[968] = ~window[28][8];
assign temp[992] = window[29][0];
assign temp[993] = window[29][1];
assign temp[994] = window[29][2];
assign temp[995] = ~window[29][3];
assign temp[996] = ~window[29][4];
assign temp[997] = window[29][5];
assign temp[998] = ~window[29][6];
assign temp[999] = ~window[29][7];
assign temp[1000] = ~window[29][8];
assign temp[1024] = ~window[30][0];
assign temp[1025] = ~window[30][1];
assign temp[1026] = ~window[30][2];
assign temp[1027] = ~window[30][3];
assign temp[1028] = ~window[30][4];
assign temp[1029] = ~window[30][5];
assign temp[1030] = ~window[30][6];
assign temp[1031] = ~window[30][7];
assign temp[1032] = ~window[30][8];
assign temp[1056] = ~window[31][0];
assign temp[1057] = ~window[31][1];
assign temp[1058] = window[31][2];
assign temp[1059] = window[31][3];
assign temp[1060] = window[31][4];
assign temp[1061] = window[31][5];
assign temp[1062] = ~window[31][6];
assign temp[1063] = window[31][7];
assign temp[1064] = ~window[31][8];
assign temp[96] = ~window[0][0];
assign temp[97] = window[0][1];
assign temp[98] = window[0][2];
assign temp[99] = window[0][3];
assign temp[100] = ~window[0][4];
assign temp[101] = window[0][5];
assign temp[102] = window[0][6];
assign temp[103] = window[0][7];
assign temp[104] = window[0][8];
assign temp[128] = window[1][0];
assign temp[129] = window[1][1];
assign temp[130] = window[1][2];
assign temp[131] = window[1][3];
assign temp[132] = ~window[1][4];
assign temp[133] = ~window[1][5];
assign temp[134] = window[1][6];
assign temp[135] = window[1][7];
assign temp[136] = ~window[1][8];
assign temp[160] = window[2][0];
assign temp[161] = window[2][1];
assign temp[162] = window[2][2];
assign temp[163] = ~window[2][3];
assign temp[164] = ~window[2][4];
assign temp[165] = ~window[2][5];
assign temp[166] = ~window[2][6];
assign temp[167] = ~window[2][7];
assign temp[168] = ~window[2][8];
assign temp[192] = ~window[3][0];
assign temp[193] = window[3][1];
assign temp[194] = window[3][2];
assign temp[195] = ~window[3][3];
assign temp[196] = ~window[3][4];
assign temp[197] = ~window[3][5];
assign temp[198] = window[3][6];
assign temp[199] = window[3][7];
assign temp[200] = window[3][8];
assign temp[224] = window[4][0];
assign temp[225] = window[4][1];
assign temp[226] = window[4][2];
assign temp[227] = window[4][3];
assign temp[228] = window[4][4];
assign temp[229] = window[4][5];
assign temp[230] = window[4][6];
assign temp[231] = window[4][7];
assign temp[232] = window[4][8];
assign temp[256] = ~window[5][0];
assign temp[257] = ~window[5][1];
assign temp[258] = ~window[5][2];
assign temp[259] = ~window[5][3];
assign temp[260] = ~window[5][4];
assign temp[261] = ~window[5][5];
assign temp[262] = window[5][6];
assign temp[263] = window[5][7];
assign temp[264] = window[5][8];
assign temp[288] = ~window[6][0];
assign temp[289] = window[6][1];
assign temp[290] = window[6][2];
assign temp[291] = ~window[6][3];
assign temp[292] = window[6][4];
assign temp[293] = window[6][5];
assign temp[294] = window[6][6];
assign temp[295] = window[6][7];
assign temp[296] = ~window[6][8];
assign temp[320] = ~window[7][0];
assign temp[321] = ~window[7][1];
assign temp[322] = ~window[7][2];
assign temp[323] = window[7][3];
assign temp[324] = window[7][4];
assign temp[325] = ~window[7][5];
assign temp[326] = window[7][6];
assign temp[327] = window[7][7];
assign temp[328] = window[7][8];
assign temp[352] = window[8][0];
assign temp[353] = window[8][1];
assign temp[354] = ~window[8][2];
assign temp[355] = window[8][3];
assign temp[356] = ~window[8][4];
assign temp[357] = ~window[8][5];
assign temp[358] = window[8][6];
assign temp[359] = window[8][7];
assign temp[360] = window[8][8];
assign temp[384] = ~window[9][0];
assign temp[385] = window[9][1];
assign temp[386] = window[9][2];
assign temp[387] = ~window[9][3];
assign temp[388] = ~window[9][4];
assign temp[389] = ~window[9][5];
assign temp[390] = window[9][6];
assign temp[391] = window[9][7];
assign temp[392] = window[9][8];
assign temp[416] = window[10][0];
assign temp[417] = ~window[10][1];
assign temp[418] = ~window[10][2];
assign temp[419] = window[10][3];
assign temp[420] = window[10][4];
assign temp[421] = window[10][5];
assign temp[422] = window[10][6];
assign temp[423] = window[10][7];
assign temp[424] = window[10][8];
assign temp[448] = window[11][0];
assign temp[449] = window[11][1];
assign temp[450] = window[11][2];
assign temp[451] = window[11][3];
assign temp[452] = window[11][4];
assign temp[453] = window[11][5];
assign temp[454] = window[11][6];
assign temp[455] = window[11][7];
assign temp[456] = window[11][8];
assign temp[480] = window[12][0];
assign temp[481] = window[12][1];
assign temp[482] = window[12][2];
assign temp[483] = ~window[12][3];
assign temp[484] = ~window[12][4];
assign temp[485] = ~window[12][5];
assign temp[486] = ~window[12][6];
assign temp[487] = window[12][7];
assign temp[488] = ~window[12][8];
assign temp[512] = ~window[13][0];
assign temp[513] = window[13][1];
assign temp[514] = ~window[13][2];
assign temp[515] = ~window[13][3];
assign temp[516] = ~window[13][4];
assign temp[517] = ~window[13][5];
assign temp[518] = ~window[13][6];
assign temp[519] = ~window[13][7];
assign temp[520] = window[13][8];
assign temp[544] = window[14][0];
assign temp[545] = ~window[14][1];
assign temp[546] = ~window[14][2];
assign temp[547] = ~window[14][3];
assign temp[548] = ~window[14][4];
assign temp[549] = ~window[14][5];
assign temp[550] = window[14][6];
assign temp[551] = window[14][7];
assign temp[552] = window[14][8];
assign temp[576] = window[15][0];
assign temp[577] = ~window[15][1];
assign temp[578] = ~window[15][2];
assign temp[579] = window[15][3];
assign temp[580] = window[15][4];
assign temp[581] = window[15][5];
assign temp[582] = window[15][6];
assign temp[583] = ~window[15][7];
assign temp[584] = window[15][8];
assign temp[608] = ~window[16][0];
assign temp[609] = ~window[16][1];
assign temp[610] = ~window[16][2];
assign temp[611] = ~window[16][3];
assign temp[612] = window[16][4];
assign temp[613] = window[16][5];
assign temp[614] = window[16][6];
assign temp[615] = window[16][7];
assign temp[616] = window[16][8];
assign temp[640] = window[17][0];
assign temp[641] = window[17][1];
assign temp[642] = window[17][2];
assign temp[643] = ~window[17][3];
assign temp[644] = ~window[17][4];
assign temp[645] = ~window[17][5];
assign temp[646] = window[17][6];
assign temp[647] = window[17][7];
assign temp[648] = ~window[17][8];
assign temp[672] = window[18][0];
assign temp[673] = ~window[18][1];
assign temp[674] = window[18][2];
assign temp[675] = ~window[18][3];
assign temp[676] = ~window[18][4];
assign temp[677] = ~window[18][5];
assign temp[678] = ~window[18][6];
assign temp[679] = window[18][7];
assign temp[680] = ~window[18][8];
assign temp[704] = window[19][0];
assign temp[705] = window[19][1];
assign temp[706] = window[19][2];
assign temp[707] = ~window[19][3];
assign temp[708] = ~window[19][4];
assign temp[709] = window[19][5];
assign temp[710] = ~window[19][6];
assign temp[711] = window[19][7];
assign temp[712] = ~window[19][8];
assign temp[736] = ~window[20][0];
assign temp[737] = window[20][1];
assign temp[738] = window[20][2];
assign temp[739] = ~window[20][3];
assign temp[740] = ~window[20][4];
assign temp[741] = ~window[20][5];
assign temp[742] = ~window[20][6];
assign temp[743] = window[20][7];
assign temp[744] = window[20][8];
assign temp[768] = ~window[21][0];
assign temp[769] = ~window[21][1];
assign temp[770] = window[21][2];
assign temp[771] = window[21][3];
assign temp[772] = ~window[21][4];
assign temp[773] = window[21][5];
assign temp[774] = window[21][6];
assign temp[775] = ~window[21][7];
assign temp[776] = ~window[21][8];
assign temp[800] = ~window[22][0];
assign temp[801] = ~window[22][1];
assign temp[802] = ~window[22][2];
assign temp[803] = window[22][3];
assign temp[804] = window[22][4];
assign temp[805] = window[22][5];
assign temp[806] = ~window[22][6];
assign temp[807] = ~window[22][7];
assign temp[808] = ~window[22][8];
assign temp[832] = ~window[23][0];
assign temp[833] = ~window[23][1];
assign temp[834] = window[23][2];
assign temp[835] = window[23][3];
assign temp[836] = ~window[23][4];
assign temp[837] = ~window[23][5];
assign temp[838] = window[23][6];
assign temp[839] = ~window[23][7];
assign temp[840] = window[23][8];
assign temp[864] = ~window[24][0];
assign temp[865] = window[24][1];
assign temp[866] = window[24][2];
assign temp[867] = ~window[24][3];
assign temp[868] = ~window[24][4];
assign temp[869] = ~window[24][5];
assign temp[870] = window[24][6];
assign temp[871] = window[24][7];
assign temp[872] = window[24][8];
assign temp[896] = ~window[25][0];
assign temp[897] = ~window[25][1];
assign temp[898] = window[25][2];
assign temp[899] = ~window[25][3];
assign temp[900] = ~window[25][4];
assign temp[901] = ~window[25][5];
assign temp[902] = window[25][6];
assign temp[903] = window[25][7];
assign temp[904] = window[25][8];
assign temp[928] = window[26][0];
assign temp[929] = ~window[26][1];
assign temp[930] = window[26][2];
assign temp[931] = window[26][3];
assign temp[932] = ~window[26][4];
assign temp[933] = ~window[26][5];
assign temp[934] = ~window[26][6];
assign temp[935] = ~window[26][7];
assign temp[936] = ~window[26][8];
assign temp[960] = window[27][0];
assign temp[961] = ~window[27][1];
assign temp[962] = ~window[27][2];
assign temp[963] = window[27][3];
assign temp[964] = window[27][4];
assign temp[965] = window[27][5];
assign temp[966] = window[27][6];
assign temp[967] = window[27][7];
assign temp[968] = window[27][8];
assign temp[992] = ~window[28][0];
assign temp[993] = window[28][1];
assign temp[994] = ~window[28][2];
assign temp[995] = window[28][3];
assign temp[996] = window[28][4];
assign temp[997] = ~window[28][5];
assign temp[998] = ~window[28][6];
assign temp[999] = ~window[28][7];
assign temp[1000] = window[28][8];
assign temp[1024] = window[29][0];
assign temp[1025] = ~window[29][1];
assign temp[1026] = ~window[29][2];
assign temp[1027] = window[29][3];
assign temp[1028] = window[29][4];
assign temp[1029] = ~window[29][5];
assign temp[1030] = ~window[29][6];
assign temp[1031] = window[29][7];
assign temp[1032] = window[29][8];
assign temp[1056] = ~window[30][0];
assign temp[1057] = ~window[30][1];
assign temp[1058] = ~window[30][2];
assign temp[1059] = ~window[30][3];
assign temp[1060] = ~window[30][4];
assign temp[1061] = ~window[30][5];
assign temp[1062] = ~window[30][6];
assign temp[1063] = ~window[30][7];
assign temp[1064] = ~window[30][8];
assign temp[1088] = window[31][0];
assign temp[1089] = window[31][1];
assign temp[1090] = window[31][2];
assign temp[1091] = ~window[31][3];
assign temp[1092] = ~window[31][4];
assign temp[1093] = ~window[31][5];
assign temp[1094] = ~window[31][6];
assign temp[1095] = window[31][7];
assign temp[1096] = window[31][8];
assign temp[128] = window[0][0];
assign temp[129] = ~window[0][1];
assign temp[130] = ~window[0][2];
assign temp[131] = ~window[0][3];
assign temp[132] = ~window[0][4];
assign temp[133] = ~window[0][5];
assign temp[134] = ~window[0][6];
assign temp[135] = ~window[0][7];
assign temp[136] = window[0][8];
assign temp[160] = window[1][0];
assign temp[161] = window[1][1];
assign temp[162] = ~window[1][2];
assign temp[163] = window[1][3];
assign temp[164] = ~window[1][4];
assign temp[165] = ~window[1][5];
assign temp[166] = window[1][6];
assign temp[167] = window[1][7];
assign temp[168] = window[1][8];
assign temp[192] = ~window[2][0];
assign temp[193] = window[2][1];
assign temp[194] = ~window[2][2];
assign temp[195] = window[2][3];
assign temp[196] = ~window[2][4];
assign temp[197] = ~window[2][5];
assign temp[198] = ~window[2][6];
assign temp[199] = window[2][7];
assign temp[200] = window[2][8];
assign temp[224] = window[3][0];
assign temp[225] = ~window[3][1];
assign temp[226] = ~window[3][2];
assign temp[227] = ~window[3][3];
assign temp[228] = ~window[3][4];
assign temp[229] = ~window[3][5];
assign temp[230] = ~window[3][6];
assign temp[231] = ~window[3][7];
assign temp[232] = window[3][8];
assign temp[256] = window[4][0];
assign temp[257] = ~window[4][1];
assign temp[258] = ~window[4][2];
assign temp[259] = ~window[4][3];
assign temp[260] = ~window[4][4];
assign temp[261] = window[4][5];
assign temp[262] = ~window[4][6];
assign temp[263] = window[4][7];
assign temp[264] = ~window[4][8];
assign temp[288] = window[5][0];
assign temp[289] = window[5][1];
assign temp[290] = ~window[5][2];
assign temp[291] = ~window[5][3];
assign temp[292] = ~window[5][4];
assign temp[293] = window[5][5];
assign temp[294] = ~window[5][6];
assign temp[295] = ~window[5][7];
assign temp[296] = window[5][8];
assign temp[320] = ~window[6][0];
assign temp[321] = ~window[6][1];
assign temp[322] = ~window[6][2];
assign temp[323] = ~window[6][3];
assign temp[324] = ~window[6][4];
assign temp[325] = window[6][5];
assign temp[326] = ~window[6][6];
assign temp[327] = window[6][7];
assign temp[328] = window[6][8];
assign temp[352] = window[7][0];
assign temp[353] = ~window[7][1];
assign temp[354] = ~window[7][2];
assign temp[355] = ~window[7][3];
assign temp[356] = ~window[7][4];
assign temp[357] = window[7][5];
assign temp[358] = ~window[7][6];
assign temp[359] = ~window[7][7];
assign temp[360] = window[7][8];
assign temp[384] = window[8][0];
assign temp[385] = ~window[8][1];
assign temp[386] = ~window[8][2];
assign temp[387] = ~window[8][3];
assign temp[388] = ~window[8][4];
assign temp[389] = window[8][5];
assign temp[390] = ~window[8][6];
assign temp[391] = window[8][7];
assign temp[392] = window[8][8];
assign temp[416] = window[9][0];
assign temp[417] = window[9][1];
assign temp[418] = ~window[9][2];
assign temp[419] = window[9][3];
assign temp[420] = ~window[9][4];
assign temp[421] = ~window[9][5];
assign temp[422] = ~window[9][6];
assign temp[423] = ~window[9][7];
assign temp[424] = ~window[9][8];
assign temp[448] = window[10][0];
assign temp[449] = window[10][1];
assign temp[450] = ~window[10][2];
assign temp[451] = ~window[10][3];
assign temp[452] = ~window[10][4];
assign temp[453] = ~window[10][5];
assign temp[454] = ~window[10][6];
assign temp[455] = ~window[10][7];
assign temp[456] = ~window[10][8];
assign temp[480] = window[11][0];
assign temp[481] = window[11][1];
assign temp[482] = window[11][2];
assign temp[483] = window[11][3];
assign temp[484] = window[11][4];
assign temp[485] = ~window[11][5];
assign temp[486] = ~window[11][6];
assign temp[487] = ~window[11][7];
assign temp[488] = ~window[11][8];
assign temp[512] = ~window[12][0];
assign temp[513] = window[12][1];
assign temp[514] = window[12][2];
assign temp[515] = window[12][3];
assign temp[516] = window[12][4];
assign temp[517] = ~window[12][5];
assign temp[518] = window[12][6];
assign temp[519] = ~window[12][7];
assign temp[520] = window[12][8];
assign temp[544] = window[13][0];
assign temp[545] = window[13][1];
assign temp[546] = window[13][2];
assign temp[547] = window[13][3];
assign temp[548] = window[13][4];
assign temp[549] = window[13][5];
assign temp[550] = window[13][6];
assign temp[551] = window[13][7];
assign temp[552] = window[13][8];
assign temp[576] = ~window[14][0];
assign temp[577] = ~window[14][1];
assign temp[578] = ~window[14][2];
assign temp[579] = ~window[14][3];
assign temp[580] = ~window[14][4];
assign temp[581] = ~window[14][5];
assign temp[582] = ~window[14][6];
assign temp[583] = ~window[14][7];
assign temp[584] = ~window[14][8];
assign temp[608] = window[15][0];
assign temp[609] = ~window[15][1];
assign temp[610] = ~window[15][2];
assign temp[611] = ~window[15][3];
assign temp[612] = ~window[15][4];
assign temp[613] = window[15][5];
assign temp[614] = ~window[15][6];
assign temp[615] = window[15][7];
assign temp[616] = ~window[15][8];
assign temp[640] = ~window[16][0];
assign temp[641] = ~window[16][1];
assign temp[642] = ~window[16][2];
assign temp[643] = ~window[16][3];
assign temp[644] = window[16][4];
assign temp[645] = ~window[16][5];
assign temp[646] = ~window[16][6];
assign temp[647] = window[16][7];
assign temp[648] = window[16][8];
assign temp[672] = window[17][0];
assign temp[673] = window[17][1];
assign temp[674] = window[17][2];
assign temp[675] = window[17][3];
assign temp[676] = ~window[17][4];
assign temp[677] = ~window[17][5];
assign temp[678] = ~window[17][6];
assign temp[679] = ~window[17][7];
assign temp[680] = window[17][8];
assign temp[704] = ~window[18][0];
assign temp[705] = window[18][1];
assign temp[706] = ~window[18][2];
assign temp[707] = window[18][3];
assign temp[708] = window[18][4];
assign temp[709] = ~window[18][5];
assign temp[710] = ~window[18][6];
assign temp[711] = window[18][7];
assign temp[712] = ~window[18][8];
assign temp[736] = ~window[19][0];
assign temp[737] = window[19][1];
assign temp[738] = window[19][2];
assign temp[739] = window[19][3];
assign temp[740] = window[19][4];
assign temp[741] = ~window[19][5];
assign temp[742] = window[19][6];
assign temp[743] = window[19][7];
assign temp[744] = ~window[19][8];
assign temp[768] = window[20][0];
assign temp[769] = window[20][1];
assign temp[770] = ~window[20][2];
assign temp[771] = ~window[20][3];
assign temp[772] = ~window[20][4];
assign temp[773] = ~window[20][5];
assign temp[774] = ~window[20][6];
assign temp[775] = ~window[20][7];
assign temp[776] = window[20][8];
assign temp[800] = window[21][0];
assign temp[801] = window[21][1];
assign temp[802] = ~window[21][2];
assign temp[803] = window[21][3];
assign temp[804] = window[21][4];
assign temp[805] = ~window[21][5];
assign temp[806] = window[21][6];
assign temp[807] = window[21][7];
assign temp[808] = window[21][8];
assign temp[832] = ~window[22][0];
assign temp[833] = ~window[22][1];
assign temp[834] = ~window[22][2];
assign temp[835] = ~window[22][3];
assign temp[836] = window[22][4];
assign temp[837] = window[22][5];
assign temp[838] = window[22][6];
assign temp[839] = window[22][7];
assign temp[840] = ~window[22][8];
assign temp[864] = window[23][0];
assign temp[865] = ~window[23][1];
assign temp[866] = ~window[23][2];
assign temp[867] = window[23][3];
assign temp[868] = window[23][4];
assign temp[869] = ~window[23][5];
assign temp[870] = ~window[23][6];
assign temp[871] = ~window[23][7];
assign temp[872] = ~window[23][8];
assign temp[896] = ~window[24][0];
assign temp[897] = window[24][1];
assign temp[898] = ~window[24][2];
assign temp[899] = ~window[24][3];
assign temp[900] = ~window[24][4];
assign temp[901] = ~window[24][5];
assign temp[902] = ~window[24][6];
assign temp[903] = ~window[24][7];
assign temp[904] = window[24][8];
assign temp[928] = ~window[25][0];
assign temp[929] = ~window[25][1];
assign temp[930] = ~window[25][2];
assign temp[931] = ~window[25][3];
assign temp[932] = window[25][4];
assign temp[933] = window[25][5];
assign temp[934] = window[25][6];
assign temp[935] = window[25][7];
assign temp[936] = window[25][8];
assign temp[960] = window[26][0];
assign temp[961] = window[26][1];
assign temp[962] = ~window[26][2];
assign temp[963] = window[26][3];
assign temp[964] = window[26][4];
assign temp[965] = window[26][5];
assign temp[966] = window[26][6];
assign temp[967] = ~window[26][7];
assign temp[968] = window[26][8];
assign temp[992] = ~window[27][0];
assign temp[993] = ~window[27][1];
assign temp[994] = ~window[27][2];
assign temp[995] = ~window[27][3];
assign temp[996] = ~window[27][4];
assign temp[997] = window[27][5];
assign temp[998] = ~window[27][6];
assign temp[999] = window[27][7];
assign temp[1000] = window[27][8];
assign temp[1024] = ~window[28][0];
assign temp[1025] = window[28][1];
assign temp[1026] = window[28][2];
assign temp[1027] = ~window[28][3];
assign temp[1028] = window[28][4];
assign temp[1029] = window[28][5];
assign temp[1030] = window[28][6];
assign temp[1031] = window[28][7];
assign temp[1032] = ~window[28][8];
assign temp[1056] = window[29][0];
assign temp[1057] = window[29][1];
assign temp[1058] = ~window[29][2];
assign temp[1059] = window[29][3];
assign temp[1060] = window[29][4];
assign temp[1061] = window[29][5];
assign temp[1062] = window[29][6];
assign temp[1063] = ~window[29][7];
assign temp[1064] = window[29][8];
assign temp[1088] = window[30][0];
assign temp[1089] = window[30][1];
assign temp[1090] = window[30][2];
assign temp[1091] = window[30][3];
assign temp[1092] = window[30][4];
assign temp[1093] = window[30][5];
assign temp[1094] = window[30][6];
assign temp[1095] = window[30][7];
assign temp[1096] = window[30][8];
assign temp[1120] = window[31][0];
assign temp[1121] = window[31][1];
assign temp[1122] = window[31][2];
assign temp[1123] = window[31][3];
assign temp[1124] = window[31][4];
assign temp[1125] = window[31][5];
assign temp[1126] = window[31][6];
assign temp[1127] = ~window[31][7];
assign temp[1128] = window[31][8];
assign temp[160] = window[0][0];
assign temp[161] = ~window[0][1];
assign temp[162] = ~window[0][2];
assign temp[163] = ~window[0][3];
assign temp[164] = ~window[0][4];
assign temp[165] = window[0][5];
assign temp[166] = ~window[0][6];
assign temp[167] = window[0][7];
assign temp[168] = window[0][8];
assign temp[192] = window[1][0];
assign temp[193] = window[1][1];
assign temp[194] = ~window[1][2];
assign temp[195] = ~window[1][3];
assign temp[196] = ~window[1][4];
assign temp[197] = ~window[1][5];
assign temp[198] = ~window[1][6];
assign temp[199] = ~window[1][7];
assign temp[200] = window[1][8];
assign temp[224] = window[2][0];
assign temp[225] = window[2][1];
assign temp[226] = ~window[2][2];
assign temp[227] = window[2][3];
assign temp[228] = ~window[2][4];
assign temp[229] = ~window[2][5];
assign temp[230] = ~window[2][6];
assign temp[231] = ~window[2][7];
assign temp[232] = window[2][8];
assign temp[256] = window[3][0];
assign temp[257] = ~window[3][1];
assign temp[258] = window[3][2];
assign temp[259] = ~window[3][3];
assign temp[260] = ~window[3][4];
assign temp[261] = window[3][5];
assign temp[262] = ~window[3][6];
assign temp[263] = window[3][7];
assign temp[264] = window[3][8];
assign temp[288] = window[4][0];
assign temp[289] = ~window[4][1];
assign temp[290] = ~window[4][2];
assign temp[291] = ~window[4][3];
assign temp[292] = ~window[4][4];
assign temp[293] = ~window[4][5];
assign temp[294] = ~window[4][6];
assign temp[295] = window[4][7];
assign temp[296] = ~window[4][8];
assign temp[320] = window[5][0];
assign temp[321] = ~window[5][1];
assign temp[322] = window[5][2];
assign temp[323] = ~window[5][3];
assign temp[324] = window[5][4];
assign temp[325] = window[5][5];
assign temp[326] = ~window[5][6];
assign temp[327] = window[5][7];
assign temp[328] = window[5][8];
assign temp[352] = window[6][0];
assign temp[353] = window[6][1];
assign temp[354] = ~window[6][2];
assign temp[355] = window[6][3];
assign temp[356] = window[6][4];
assign temp[357] = ~window[6][5];
assign temp[358] = window[6][6];
assign temp[359] = ~window[6][7];
assign temp[360] = ~window[6][8];
assign temp[384] = ~window[7][0];
assign temp[385] = ~window[7][1];
assign temp[386] = window[7][2];
assign temp[387] = ~window[7][3];
assign temp[388] = window[7][4];
assign temp[389] = window[7][5];
assign temp[390] = ~window[7][6];
assign temp[391] = window[7][7];
assign temp[392] = window[7][8];
assign temp[416] = ~window[8][0];
assign temp[417] = ~window[8][1];
assign temp[418] = ~window[8][2];
assign temp[419] = ~window[8][3];
assign temp[420] = ~window[8][4];
assign temp[421] = window[8][5];
assign temp[422] = window[8][6];
assign temp[423] = window[8][7];
assign temp[424] = window[8][8];
assign temp[448] = window[9][0];
assign temp[449] = ~window[9][1];
assign temp[450] = ~window[9][2];
assign temp[451] = ~window[9][3];
assign temp[452] = ~window[9][4];
assign temp[453] = window[9][5];
assign temp[454] = ~window[9][6];
assign temp[455] = window[9][7];
assign temp[456] = window[9][8];
assign temp[480] = window[10][0];
assign temp[481] = ~window[10][1];
assign temp[482] = ~window[10][2];
assign temp[483] = ~window[10][3];
assign temp[484] = ~window[10][4];
assign temp[485] = window[10][5];
assign temp[486] = ~window[10][6];
assign temp[487] = ~window[10][7];
assign temp[488] = window[10][8];
assign temp[512] = ~window[11][0];
assign temp[513] = ~window[11][1];
assign temp[514] = window[11][2];
assign temp[515] = window[11][3];
assign temp[516] = ~window[11][4];
assign temp[517] = ~window[11][5];
assign temp[518] = ~window[11][6];
assign temp[519] = window[11][7];
assign temp[520] = window[11][8];
assign temp[544] = ~window[12][0];
assign temp[545] = ~window[12][1];
assign temp[546] = ~window[12][2];
assign temp[547] = window[12][3];
assign temp[548] = ~window[12][4];
assign temp[549] = window[12][5];
assign temp[550] = window[12][6];
assign temp[551] = ~window[12][7];
assign temp[552] = window[12][8];
assign temp[576] = ~window[13][0];
assign temp[577] = ~window[13][1];
assign temp[578] = ~window[13][2];
assign temp[579] = window[13][3];
assign temp[580] = window[13][4];
assign temp[581] = window[13][5];
assign temp[582] = window[13][6];
assign temp[583] = window[13][7];
assign temp[584] = window[13][8];
assign temp[608] = ~window[14][0];
assign temp[609] = ~window[14][1];
assign temp[610] = ~window[14][2];
assign temp[611] = ~window[14][3];
assign temp[612] = ~window[14][4];
assign temp[613] = window[14][5];
assign temp[614] = window[14][6];
assign temp[615] = window[14][7];
assign temp[616] = window[14][8];
assign temp[640] = ~window[15][0];
assign temp[641] = ~window[15][1];
assign temp[642] = window[15][2];
assign temp[643] = window[15][3];
assign temp[644] = window[15][4];
assign temp[645] = ~window[15][5];
assign temp[646] = window[15][6];
assign temp[647] = ~window[15][7];
assign temp[648] = ~window[15][8];
assign temp[672] = ~window[16][0];
assign temp[673] = window[16][1];
assign temp[674] = window[16][2];
assign temp[675] = ~window[16][3];
assign temp[676] = window[16][4];
assign temp[677] = window[16][5];
assign temp[678] = window[16][6];
assign temp[679] = window[16][7];
assign temp[680] = window[16][8];
assign temp[704] = window[17][0];
assign temp[705] = window[17][1];
assign temp[706] = ~window[17][2];
assign temp[707] = ~window[17][3];
assign temp[708] = ~window[17][4];
assign temp[709] = ~window[17][5];
assign temp[710] = ~window[17][6];
assign temp[711] = window[17][7];
assign temp[712] = window[17][8];
assign temp[736] = window[18][0];
assign temp[737] = window[18][1];
assign temp[738] = window[18][2];
assign temp[739] = window[18][3];
assign temp[740] = ~window[18][4];
assign temp[741] = window[18][5];
assign temp[742] = ~window[18][6];
assign temp[743] = ~window[18][7];
assign temp[744] = ~window[18][8];
assign temp[768] = window[19][0];
assign temp[769] = window[19][1];
assign temp[770] = ~window[19][2];
assign temp[771] = ~window[19][3];
assign temp[772] = ~window[19][4];
assign temp[773] = window[19][5];
assign temp[774] = ~window[19][6];
assign temp[775] = window[19][7];
assign temp[776] = ~window[19][8];
assign temp[800] = window[20][0];
assign temp[801] = ~window[20][1];
assign temp[802] = window[20][2];
assign temp[803] = ~window[20][3];
assign temp[804] = ~window[20][4];
assign temp[805] = window[20][5];
assign temp[806] = ~window[20][6];
assign temp[807] = window[20][7];
assign temp[808] = window[20][8];
assign temp[832] = window[21][0];
assign temp[833] = ~window[21][1];
assign temp[834] = ~window[21][2];
assign temp[835] = ~window[21][3];
assign temp[836] = ~window[21][4];
assign temp[837] = ~window[21][5];
assign temp[838] = ~window[21][6];
assign temp[839] = ~window[21][7];
assign temp[840] = ~window[21][8];
assign temp[864] = window[22][0];
assign temp[865] = window[22][1];
assign temp[866] = ~window[22][2];
assign temp[867] = window[22][3];
assign temp[868] = window[22][4];
assign temp[869] = ~window[22][5];
assign temp[870] = window[22][6];
assign temp[871] = ~window[22][7];
assign temp[872] = ~window[22][8];
assign temp[896] = ~window[23][0];
assign temp[897] = ~window[23][1];
assign temp[898] = window[23][2];
assign temp[899] = window[23][3];
assign temp[900] = window[23][4];
assign temp[901] = window[23][5];
assign temp[902] = ~window[23][6];
assign temp[903] = window[23][7];
assign temp[904] = window[23][8];
assign temp[928] = window[24][0];
assign temp[929] = ~window[24][1];
assign temp[930] = ~window[24][2];
assign temp[931] = window[24][3];
assign temp[932] = ~window[24][4];
assign temp[933] = window[24][5];
assign temp[934] = ~window[24][6];
assign temp[935] = ~window[24][7];
assign temp[936] = window[24][8];
assign temp[960] = ~window[25][0];
assign temp[961] = ~window[25][1];
assign temp[962] = ~window[25][2];
assign temp[963] = ~window[25][3];
assign temp[964] = window[25][4];
assign temp[965] = window[25][5];
assign temp[966] = window[25][6];
assign temp[967] = window[25][7];
assign temp[968] = window[25][8];
assign temp[992] = window[26][0];
assign temp[993] = ~window[26][1];
assign temp[994] = ~window[26][2];
assign temp[995] = window[26][3];
assign temp[996] = ~window[26][4];
assign temp[997] = ~window[26][5];
assign temp[998] = ~window[26][6];
assign temp[999] = window[26][7];
assign temp[1000] = ~window[26][8];
assign temp[1024] = ~window[27][0];
assign temp[1025] = ~window[27][1];
assign temp[1026] = ~window[27][2];
assign temp[1027] = ~window[27][3];
assign temp[1028] = window[27][4];
assign temp[1029] = window[27][5];
assign temp[1030] = window[27][6];
assign temp[1031] = window[27][7];
assign temp[1032] = ~window[27][8];
assign temp[1056] = ~window[28][0];
assign temp[1057] = ~window[28][1];
assign temp[1058] = ~window[28][2];
assign temp[1059] = window[28][3];
assign temp[1060] = window[28][4];
assign temp[1061] = window[28][5];
assign temp[1062] = window[28][6];
assign temp[1063] = window[28][7];
assign temp[1064] = window[28][8];
assign temp[1088] = ~window[29][0];
assign temp[1089] = ~window[29][1];
assign temp[1090] = ~window[29][2];
assign temp[1091] = window[29][3];
assign temp[1092] = ~window[29][4];
assign temp[1093] = ~window[29][5];
assign temp[1094] = window[29][6];
assign temp[1095] = window[29][7];
assign temp[1096] = window[29][8];
assign temp[1120] = window[30][0];
assign temp[1121] = ~window[30][1];
assign temp[1122] = window[30][2];
assign temp[1123] = window[30][3];
assign temp[1124] = window[30][4];
assign temp[1125] = window[30][5];
assign temp[1126] = window[30][6];
assign temp[1127] = window[30][7];
assign temp[1128] = window[30][8];
assign temp[1152] = window[31][0];
assign temp[1153] = window[31][1];
assign temp[1154] = ~window[31][2];
assign temp[1155] = window[31][3];
assign temp[1156] = ~window[31][4];
assign temp[1157] = window[31][5];
assign temp[1158] = ~window[31][6];
assign temp[1159] = ~window[31][7];
assign temp[1160] = window[31][8];
assign temp[192] = window[0][0];
assign temp[193] = window[0][1];
assign temp[194] = window[0][2];
assign temp[195] = ~window[0][3];
assign temp[196] = ~window[0][4];
assign temp[197] = window[0][5];
assign temp[198] = window[0][6];
assign temp[199] = window[0][7];
assign temp[200] = window[0][8];
assign temp[224] = window[1][0];
assign temp[225] = window[1][1];
assign temp[226] = ~window[1][2];
assign temp[227] = window[1][3];
assign temp[228] = ~window[1][4];
assign temp[229] = window[1][5];
assign temp[230] = window[1][6];
assign temp[231] = window[1][7];
assign temp[232] = window[1][8];
assign temp[256] = window[2][0];
assign temp[257] = ~window[2][1];
assign temp[258] = window[2][2];
assign temp[259] = window[2][3];
assign temp[260] = window[2][4];
assign temp[261] = window[2][5];
assign temp[262] = window[2][6];
assign temp[263] = window[2][7];
assign temp[264] = window[2][8];
assign temp[288] = window[3][0];
assign temp[289] = ~window[3][1];
assign temp[290] = window[3][2];
assign temp[291] = window[3][3];
assign temp[292] = window[3][4];
assign temp[293] = window[3][5];
assign temp[294] = ~window[3][6];
assign temp[295] = ~window[3][7];
assign temp[296] = ~window[3][8];
assign temp[320] = window[4][0];
assign temp[321] = window[4][1];
assign temp[322] = window[4][2];
assign temp[323] = ~window[4][3];
assign temp[324] = ~window[4][4];
assign temp[325] = ~window[4][5];
assign temp[326] = ~window[4][6];
assign temp[327] = ~window[4][7];
assign temp[328] = ~window[4][8];
assign temp[352] = window[5][0];
assign temp[353] = window[5][1];
assign temp[354] = window[5][2];
assign temp[355] = ~window[5][3];
assign temp[356] = window[5][4];
assign temp[357] = window[5][5];
assign temp[358] = ~window[5][6];
assign temp[359] = ~window[5][7];
assign temp[360] = ~window[5][8];
assign temp[384] = ~window[6][0];
assign temp[385] = ~window[6][1];
assign temp[386] = ~window[6][2];
assign temp[387] = window[6][3];
assign temp[388] = ~window[6][4];
assign temp[389] = window[6][5];
assign temp[390] = window[6][6];
assign temp[391] = window[6][7];
assign temp[392] = window[6][8];
assign temp[416] = window[7][0];
assign temp[417] = ~window[7][1];
assign temp[418] = window[7][2];
assign temp[419] = ~window[7][3];
assign temp[420] = ~window[7][4];
assign temp[421] = ~window[7][5];
assign temp[422] = ~window[7][6];
assign temp[423] = ~window[7][7];
assign temp[424] = ~window[7][8];
assign temp[448] = window[8][0];
assign temp[449] = window[8][1];
assign temp[450] = window[8][2];
assign temp[451] = window[8][3];
assign temp[452] = ~window[8][4];
assign temp[453] = window[8][5];
assign temp[454] = window[8][6];
assign temp[455] = window[8][7];
assign temp[456] = window[8][8];
assign temp[480] = ~window[9][0];
assign temp[481] = ~window[9][1];
assign temp[482] = window[9][2];
assign temp[483] = window[9][3];
assign temp[484] = window[9][4];
assign temp[485] = window[9][5];
assign temp[486] = ~window[9][6];
assign temp[487] = ~window[9][7];
assign temp[488] = ~window[9][8];
assign temp[512] = window[10][0];
assign temp[513] = ~window[10][1];
assign temp[514] = ~window[10][2];
assign temp[515] = ~window[10][3];
assign temp[516] = ~window[10][4];
assign temp[517] = ~window[10][5];
assign temp[518] = ~window[10][6];
assign temp[519] = ~window[10][7];
assign temp[520] = ~window[10][8];
assign temp[544] = window[11][0];
assign temp[545] = ~window[11][1];
assign temp[546] = ~window[11][2];
assign temp[547] = ~window[11][3];
assign temp[548] = window[11][4];
assign temp[549] = ~window[11][5];
assign temp[550] = ~window[11][6];
assign temp[551] = ~window[11][7];
assign temp[552] = ~window[11][8];
assign temp[576] = ~window[12][0];
assign temp[577] = window[12][1];
assign temp[578] = ~window[12][2];
assign temp[579] = window[12][3];
assign temp[580] = ~window[12][4];
assign temp[581] = window[12][5];
assign temp[582] = window[12][6];
assign temp[583] = window[12][7];
assign temp[584] = window[12][8];
assign temp[608] = ~window[13][0];
assign temp[609] = window[13][1];
assign temp[610] = ~window[13][2];
assign temp[611] = window[13][3];
assign temp[612] = window[13][4];
assign temp[613] = window[13][5];
assign temp[614] = ~window[13][6];
assign temp[615] = ~window[13][7];
assign temp[616] = ~window[13][8];
assign temp[640] = ~window[14][0];
assign temp[641] = window[14][1];
assign temp[642] = window[14][2];
assign temp[643] = window[14][3];
assign temp[644] = window[14][4];
assign temp[645] = ~window[14][5];
assign temp[646] = window[14][6];
assign temp[647] = ~window[14][7];
assign temp[648] = ~window[14][8];
assign temp[672] = window[15][0];
assign temp[673] = window[15][1];
assign temp[674] = ~window[15][2];
assign temp[675] = window[15][3];
assign temp[676] = ~window[15][4];
assign temp[677] = ~window[15][5];
assign temp[678] = window[15][6];
assign temp[679] = window[15][7];
assign temp[680] = ~window[15][8];
assign temp[704] = ~window[16][0];
assign temp[705] = window[16][1];
assign temp[706] = window[16][2];
assign temp[707] = ~window[16][3];
assign temp[708] = ~window[16][4];
assign temp[709] = window[16][5];
assign temp[710] = ~window[16][6];
assign temp[711] = ~window[16][7];
assign temp[712] = ~window[16][8];
assign temp[736] = window[17][0];
assign temp[737] = window[17][1];
assign temp[738] = window[17][2];
assign temp[739] = window[17][3];
assign temp[740] = window[17][4];
assign temp[741] = window[17][5];
assign temp[742] = ~window[17][6];
assign temp[743] = window[17][7];
assign temp[744] = window[17][8];
assign temp[768] = window[18][0];
assign temp[769] = window[18][1];
assign temp[770] = window[18][2];
assign temp[771] = ~window[18][3];
assign temp[772] = window[18][4];
assign temp[773] = window[18][5];
assign temp[774] = ~window[18][6];
assign temp[775] = ~window[18][7];
assign temp[776] = ~window[18][8];
assign temp[800] = window[19][0];
assign temp[801] = window[19][1];
assign temp[802] = ~window[19][2];
assign temp[803] = window[19][3];
assign temp[804] = window[19][4];
assign temp[805] = ~window[19][5];
assign temp[806] = window[19][6];
assign temp[807] = ~window[19][7];
assign temp[808] = ~window[19][8];
assign temp[832] = window[20][0];
assign temp[833] = ~window[20][1];
assign temp[834] = window[20][2];
assign temp[835] = window[20][3];
assign temp[836] = window[20][4];
assign temp[837] = window[20][5];
assign temp[838] = ~window[20][6];
assign temp[839] = ~window[20][7];
assign temp[840] = ~window[20][8];
assign temp[864] = window[21][0];
assign temp[865] = window[21][1];
assign temp[866] = ~window[21][2];
assign temp[867] = ~window[21][3];
assign temp[868] = ~window[21][4];
assign temp[869] = ~window[21][5];
assign temp[870] = ~window[21][6];
assign temp[871] = ~window[21][7];
assign temp[872] = ~window[21][8];
assign temp[896] = ~window[22][0];
assign temp[897] = window[22][1];
assign temp[898] = ~window[22][2];
assign temp[899] = window[22][3];
assign temp[900] = ~window[22][4];
assign temp[901] = ~window[22][5];
assign temp[902] = window[22][6];
assign temp[903] = window[22][7];
assign temp[904] = window[22][8];
assign temp[928] = ~window[23][0];
assign temp[929] = window[23][1];
assign temp[930] = window[23][2];
assign temp[931] = ~window[23][3];
assign temp[932] = ~window[23][4];
assign temp[933] = window[23][5];
assign temp[934] = ~window[23][6];
assign temp[935] = ~window[23][7];
assign temp[936] = ~window[23][8];
assign temp[960] = window[24][0];
assign temp[961] = ~window[24][1];
assign temp[962] = window[24][2];
assign temp[963] = window[24][3];
assign temp[964] = window[24][4];
assign temp[965] = window[24][5];
assign temp[966] = ~window[24][6];
assign temp[967] = window[24][7];
assign temp[968] = window[24][8];
assign temp[992] = ~window[25][0];
assign temp[993] = window[25][1];
assign temp[994] = window[25][2];
assign temp[995] = window[25][3];
assign temp[996] = window[25][4];
assign temp[997] = window[25][5];
assign temp[998] = ~window[25][6];
assign temp[999] = ~window[25][7];
assign temp[1000] = window[25][8];
assign temp[1024] = window[26][0];
assign temp[1025] = window[26][1];
assign temp[1026] = ~window[26][2];
assign temp[1027] = window[26][3];
assign temp[1028] = ~window[26][4];
assign temp[1029] = ~window[26][5];
assign temp[1030] = window[26][6];
assign temp[1031] = window[26][7];
assign temp[1032] = window[26][8];
assign temp[1056] = window[27][0];
assign temp[1057] = window[27][1];
assign temp[1058] = ~window[27][2];
assign temp[1059] = ~window[27][3];
assign temp[1060] = ~window[27][4];
assign temp[1061] = ~window[27][5];
assign temp[1062] = ~window[27][6];
assign temp[1063] = ~window[27][7];
assign temp[1064] = ~window[27][8];
assign temp[1088] = ~window[28][0];
assign temp[1089] = ~window[28][1];
assign temp[1090] = window[28][2];
assign temp[1091] = ~window[28][3];
assign temp[1092] = ~window[28][4];
assign temp[1093] = ~window[28][5];
assign temp[1094] = ~window[28][6];
assign temp[1095] = ~window[28][7];
assign temp[1096] = ~window[28][8];
assign temp[1120] = ~window[29][0];
assign temp[1121] = window[29][1];
assign temp[1122] = ~window[29][2];
assign temp[1123] = ~window[29][3];
assign temp[1124] = ~window[29][4];
assign temp[1125] = ~window[29][5];
assign temp[1126] = ~window[29][6];
assign temp[1127] = window[29][7];
assign temp[1128] = ~window[29][8];
assign temp[1152] = ~window[30][0];
assign temp[1153] = window[30][1];
assign temp[1154] = window[30][2];
assign temp[1155] = ~window[30][3];
assign temp[1156] = window[30][4];
assign temp[1157] = ~window[30][5];
assign temp[1158] = ~window[30][6];
assign temp[1159] = window[30][7];
assign temp[1160] = ~window[30][8];
assign temp[1184] = ~window[31][0];
assign temp[1185] = window[31][1];
assign temp[1186] = window[31][2];
assign temp[1187] = window[31][3];
assign temp[1188] = window[31][4];
assign temp[1189] = window[31][5];
assign temp[1190] = ~window[31][6];
assign temp[1191] = window[31][7];
assign temp[1192] = window[31][8];
assign temp[224] = ~window[0][0];
assign temp[225] = window[0][1];
assign temp[226] = window[0][2];
assign temp[227] = ~window[0][3];
assign temp[228] = window[0][4];
assign temp[229] = window[0][5];
assign temp[230] = ~window[0][6];
assign temp[231] = window[0][7];
assign temp[232] = window[0][8];
assign temp[256] = ~window[1][0];
assign temp[257] = ~window[1][1];
assign temp[258] = window[1][2];
assign temp[259] = window[1][3];
assign temp[260] = window[1][4];
assign temp[261] = ~window[1][5];
assign temp[262] = ~window[1][6];
assign temp[263] = ~window[1][7];
assign temp[264] = ~window[1][8];
assign temp[288] = window[2][0];
assign temp[289] = ~window[2][1];
assign temp[290] = window[2][2];
assign temp[291] = window[2][3];
assign temp[292] = window[2][4];
assign temp[293] = window[2][5];
assign temp[294] = ~window[2][6];
assign temp[295] = window[2][7];
assign temp[296] = ~window[2][8];
assign temp[320] = window[3][0];
assign temp[321] = window[3][1];
assign temp[322] = window[3][2];
assign temp[323] = window[3][3];
assign temp[324] = ~window[3][4];
assign temp[325] = window[3][5];
assign temp[326] = ~window[3][6];
assign temp[327] = ~window[3][7];
assign temp[328] = ~window[3][8];
assign temp[352] = window[4][0];
assign temp[353] = window[4][1];
assign temp[354] = window[4][2];
assign temp[355] = ~window[4][3];
assign temp[356] = ~window[4][4];
assign temp[357] = ~window[4][5];
assign temp[358] = ~window[4][6];
assign temp[359] = window[4][7];
assign temp[360] = window[4][8];
assign temp[384] = ~window[5][0];
assign temp[385] = window[5][1];
assign temp[386] = window[5][2];
assign temp[387] = ~window[5][3];
assign temp[388] = ~window[5][4];
assign temp[389] = ~window[5][5];
assign temp[390] = ~window[5][6];
assign temp[391] = ~window[5][7];
assign temp[392] = window[5][8];
assign temp[416] = ~window[6][0];
assign temp[417] = window[6][1];
assign temp[418] = ~window[6][2];
assign temp[419] = ~window[6][3];
assign temp[420] = window[6][4];
assign temp[421] = window[6][5];
assign temp[422] = window[6][6];
assign temp[423] = window[6][7];
assign temp[424] = window[6][8];
assign temp[448] = window[7][0];
assign temp[449] = window[7][1];
assign temp[450] = window[7][2];
assign temp[451] = window[7][3];
assign temp[452] = ~window[7][4];
assign temp[453] = ~window[7][5];
assign temp[454] = ~window[7][6];
assign temp[455] = window[7][7];
assign temp[456] = window[7][8];
assign temp[480] = ~window[8][0];
assign temp[481] = window[8][1];
assign temp[482] = window[8][2];
assign temp[483] = ~window[8][3];
assign temp[484] = window[8][4];
assign temp[485] = ~window[8][5];
assign temp[486] = window[8][6];
assign temp[487] = window[8][7];
assign temp[488] = window[8][8];
assign temp[512] = ~window[9][0];
assign temp[513] = window[9][1];
assign temp[514] = window[9][2];
assign temp[515] = window[9][3];
assign temp[516] = window[9][4];
assign temp[517] = window[9][5];
assign temp[518] = ~window[9][6];
assign temp[519] = ~window[9][7];
assign temp[520] = ~window[9][8];
assign temp[544] = window[10][0];
assign temp[545] = window[10][1];
assign temp[546] = window[10][2];
assign temp[547] = window[10][3];
assign temp[548] = window[10][4];
assign temp[549] = ~window[10][5];
assign temp[550] = ~window[10][6];
assign temp[551] = ~window[10][7];
assign temp[552] = window[10][8];
assign temp[576] = window[11][0];
assign temp[577] = window[11][1];
assign temp[578] = ~window[11][2];
assign temp[579] = ~window[11][3];
assign temp[580] = ~window[11][4];
assign temp[581] = ~window[11][5];
assign temp[582] = window[11][6];
assign temp[583] = window[11][7];
assign temp[584] = window[11][8];
assign temp[608] = ~window[12][0];
assign temp[609] = ~window[12][1];
assign temp[610] = ~window[12][2];
assign temp[611] = window[12][3];
assign temp[612] = window[12][4];
assign temp[613] = window[12][5];
assign temp[614] = window[12][6];
assign temp[615] = window[12][7];
assign temp[616] = ~window[12][8];
assign temp[640] = window[13][0];
assign temp[641] = ~window[13][1];
assign temp[642] = ~window[13][2];
assign temp[643] = ~window[13][3];
assign temp[644] = window[13][4];
assign temp[645] = window[13][5];
assign temp[646] = window[13][6];
assign temp[647] = window[13][7];
assign temp[648] = window[13][8];
assign temp[672] = window[14][0];
assign temp[673] = window[14][1];
assign temp[674] = ~window[14][2];
assign temp[675] = ~window[14][3];
assign temp[676] = ~window[14][4];
assign temp[677] = ~window[14][5];
assign temp[678] = window[14][6];
assign temp[679] = window[14][7];
assign temp[680] = window[14][8];
assign temp[704] = ~window[15][0];
assign temp[705] = ~window[15][1];
assign temp[706] = ~window[15][2];
assign temp[707] = ~window[15][3];
assign temp[708] = ~window[15][4];
assign temp[709] = ~window[15][5];
assign temp[710] = window[15][6];
assign temp[711] = window[15][7];
assign temp[712] = window[15][8];
assign temp[736] = window[16][0];
assign temp[737] = window[16][1];
assign temp[738] = window[16][2];
assign temp[739] = ~window[16][3];
assign temp[740] = ~window[16][4];
assign temp[741] = ~window[16][5];
assign temp[742] = window[16][6];
assign temp[743] = window[16][7];
assign temp[744] = window[16][8];
assign temp[768] = ~window[17][0];
assign temp[769] = ~window[17][1];
assign temp[770] = ~window[17][2];
assign temp[771] = window[17][3];
assign temp[772] = window[17][4];
assign temp[773] = window[17][5];
assign temp[774] = ~window[17][6];
assign temp[775] = ~window[17][7];
assign temp[776] = ~window[17][8];
assign temp[800] = ~window[18][0];
assign temp[801] = window[18][1];
assign temp[802] = window[18][2];
assign temp[803] = window[18][3];
assign temp[804] = ~window[18][4];
assign temp[805] = ~window[18][5];
assign temp[806] = ~window[18][6];
assign temp[807] = ~window[18][7];
assign temp[808] = ~window[18][8];
assign temp[832] = ~window[19][0];
assign temp[833] = ~window[19][1];
assign temp[834] = window[19][2];
assign temp[835] = window[19][3];
assign temp[836] = window[19][4];
assign temp[837] = window[19][5];
assign temp[838] = ~window[19][6];
assign temp[839] = ~window[19][7];
assign temp[840] = ~window[19][8];
assign temp[864] = ~window[20][0];
assign temp[865] = window[20][1];
assign temp[866] = window[20][2];
assign temp[867] = window[20][3];
assign temp[868] = window[20][4];
assign temp[869] = window[20][5];
assign temp[870] = ~window[20][6];
assign temp[871] = ~window[20][7];
assign temp[872] = ~window[20][8];
assign temp[896] = ~window[21][0];
assign temp[897] = ~window[21][1];
assign temp[898] = ~window[21][2];
assign temp[899] = window[21][3];
assign temp[900] = ~window[21][4];
assign temp[901] = ~window[21][5];
assign temp[902] = ~window[21][6];
assign temp[903] = ~window[21][7];
assign temp[904] = ~window[21][8];
assign temp[928] = window[22][0];
assign temp[929] = window[22][1];
assign temp[930] = window[22][2];
assign temp[931] = ~window[22][3];
assign temp[932] = ~window[22][4];
assign temp[933] = ~window[22][5];
assign temp[934] = window[22][6];
assign temp[935] = window[22][7];
assign temp[936] = window[22][8];
assign temp[960] = ~window[23][0];
assign temp[961] = ~window[23][1];
assign temp[962] = window[23][2];
assign temp[963] = ~window[23][3];
assign temp[964] = window[23][4];
assign temp[965] = ~window[23][5];
assign temp[966] = ~window[23][6];
assign temp[967] = ~window[23][7];
assign temp[968] = ~window[23][8];
assign temp[992] = window[24][0];
assign temp[993] = ~window[24][1];
assign temp[994] = window[24][2];
assign temp[995] = window[24][3];
assign temp[996] = window[24][4];
assign temp[997] = window[24][5];
assign temp[998] = ~window[24][6];
assign temp[999] = ~window[24][7];
assign temp[1000] = ~window[24][8];
assign temp[1024] = window[25][0];
assign temp[1025] = window[25][1];
assign temp[1026] = ~window[25][2];
assign temp[1027] = ~window[25][3];
assign temp[1028] = ~window[25][4];
assign temp[1029] = ~window[25][5];
assign temp[1030] = ~window[25][6];
assign temp[1031] = window[25][7];
assign temp[1032] = ~window[25][8];
assign temp[1056] = ~window[26][0];
assign temp[1057] = ~window[26][1];
assign temp[1058] = ~window[26][2];
assign temp[1059] = ~window[26][3];
assign temp[1060] = window[26][4];
assign temp[1061] = window[26][5];
assign temp[1062] = window[26][6];
assign temp[1063] = window[26][7];
assign temp[1064] = window[26][8];
assign temp[1088] = window[27][0];
assign temp[1089] = window[27][1];
assign temp[1090] = ~window[27][2];
assign temp[1091] = ~window[27][3];
assign temp[1092] = ~window[27][4];
assign temp[1093] = ~window[27][5];
assign temp[1094] = window[27][6];
assign temp[1095] = window[27][7];
assign temp[1096] = window[27][8];
assign temp[1120] = window[28][0];
assign temp[1121] = window[28][1];
assign temp[1122] = window[28][2];
assign temp[1123] = window[28][3];
assign temp[1124] = ~window[28][4];
assign temp[1125] = ~window[28][5];
assign temp[1126] = window[28][6];
assign temp[1127] = window[28][7];
assign temp[1128] = window[28][8];
assign temp[1152] = window[29][0];
assign temp[1153] = ~window[29][1];
assign temp[1154] = window[29][2];
assign temp[1155] = ~window[29][3];
assign temp[1156] = ~window[29][4];
assign temp[1157] = ~window[29][5];
assign temp[1158] = window[29][6];
assign temp[1159] = window[29][7];
assign temp[1160] = window[29][8];
assign temp[1184] = ~window[30][0];
assign temp[1185] = ~window[30][1];
assign temp[1186] = ~window[30][2];
assign temp[1187] = ~window[30][3];
assign temp[1188] = ~window[30][4];
assign temp[1189] = ~window[30][5];
assign temp[1190] = ~window[30][6];
assign temp[1191] = window[30][7];
assign temp[1192] = window[30][8];
assign temp[1216] = window[31][0];
assign temp[1217] = ~window[31][1];
assign temp[1218] = window[31][2];
assign temp[1219] = window[31][3];
assign temp[1220] = window[31][4];
assign temp[1221] = window[31][5];
assign temp[1222] = ~window[31][6];
assign temp[1223] = window[31][7];
assign temp[1224] = ~window[31][8];
assign temp[256] = window[0][0];
assign temp[257] = ~window[0][1];
assign temp[258] = ~window[0][2];
assign temp[259] = ~window[0][3];
assign temp[260] = ~window[0][4];
assign temp[261] = ~window[0][5];
assign temp[262] = window[0][6];
assign temp[263] = ~window[0][7];
assign temp[264] = ~window[0][8];
assign temp[288] = window[1][0];
assign temp[289] = window[1][1];
assign temp[290] = ~window[1][2];
assign temp[291] = window[1][3];
assign temp[292] = window[1][4];
assign temp[293] = ~window[1][5];
assign temp[294] = window[1][6];
assign temp[295] = ~window[1][7];
assign temp[296] = ~window[1][8];
assign temp[320] = window[2][0];
assign temp[321] = window[2][1];
assign temp[322] = window[2][2];
assign temp[323] = window[2][3];
assign temp[324] = ~window[2][4];
assign temp[325] = ~window[2][5];
assign temp[326] = window[2][6];
assign temp[327] = window[2][7];
assign temp[328] = window[2][8];
assign temp[352] = ~window[3][0];
assign temp[353] = ~window[3][1];
assign temp[354] = ~window[3][2];
assign temp[355] = window[3][3];
assign temp[356] = ~window[3][4];
assign temp[357] = ~window[3][5];
assign temp[358] = window[3][6];
assign temp[359] = window[3][7];
assign temp[360] = window[3][8];
assign temp[384] = window[4][0];
assign temp[385] = window[4][1];
assign temp[386] = ~window[4][2];
assign temp[387] = window[4][3];
assign temp[388] = window[4][4];
assign temp[389] = window[4][5];
assign temp[390] = window[4][6];
assign temp[391] = window[4][7];
assign temp[392] = window[4][8];
assign temp[416] = window[5][0];
assign temp[417] = ~window[5][1];
assign temp[418] = ~window[5][2];
assign temp[419] = window[5][3];
assign temp[420] = ~window[5][4];
assign temp[421] = ~window[5][5];
assign temp[422] = window[5][6];
assign temp[423] = window[5][7];
assign temp[424] = ~window[5][8];
assign temp[448] = window[6][0];
assign temp[449] = window[6][1];
assign temp[450] = ~window[6][2];
assign temp[451] = ~window[6][3];
assign temp[452] = window[6][4];
assign temp[453] = window[6][5];
assign temp[454] = ~window[6][6];
assign temp[455] = ~window[6][7];
assign temp[456] = ~window[6][8];
assign temp[480] = window[7][0];
assign temp[481] = ~window[7][1];
assign temp[482] = ~window[7][2];
assign temp[483] = window[7][3];
assign temp[484] = ~window[7][4];
assign temp[485] = ~window[7][5];
assign temp[486] = window[7][6];
assign temp[487] = window[7][7];
assign temp[488] = window[7][8];
assign temp[512] = window[8][0];
assign temp[513] = ~window[8][1];
assign temp[514] = ~window[8][2];
assign temp[515] = window[8][3];
assign temp[516] = ~window[8][4];
assign temp[517] = ~window[8][5];
assign temp[518] = window[8][6];
assign temp[519] = window[8][7];
assign temp[520] = window[8][8];
assign temp[544] = window[9][0];
assign temp[545] = window[9][1];
assign temp[546] = ~window[9][2];
assign temp[547] = window[9][3];
assign temp[548] = ~window[9][4];
assign temp[549] = ~window[9][5];
assign temp[550] = window[9][6];
assign temp[551] = window[9][7];
assign temp[552] = window[9][8];
assign temp[576] = window[10][0];
assign temp[577] = window[10][1];
assign temp[578] = ~window[10][2];
assign temp[579] = window[10][3];
assign temp[580] = window[10][4];
assign temp[581] = window[10][5];
assign temp[582] = window[10][6];
assign temp[583] = window[10][7];
assign temp[584] = window[10][8];
assign temp[608] = window[11][0];
assign temp[609] = window[11][1];
assign temp[610] = ~window[11][2];
assign temp[611] = window[11][3];
assign temp[612] = window[11][4];
assign temp[613] = window[11][5];
assign temp[614] = window[11][6];
assign temp[615] = window[11][7];
assign temp[616] = window[11][8];
assign temp[640] = window[12][0];
assign temp[641] = ~window[12][1];
assign temp[642] = ~window[12][2];
assign temp[643] = window[12][3];
assign temp[644] = window[12][4];
assign temp[645] = window[12][5];
assign temp[646] = window[12][6];
assign temp[647] = ~window[12][7];
assign temp[648] = ~window[12][8];
assign temp[672] = window[13][0];
assign temp[673] = window[13][1];
assign temp[674] = ~window[13][2];
assign temp[675] = window[13][3];
assign temp[676] = window[13][4];
assign temp[677] = window[13][5];
assign temp[678] = window[13][6];
assign temp[679] = ~window[13][7];
assign temp[680] = window[13][8];
assign temp[704] = ~window[14][0];
assign temp[705] = ~window[14][1];
assign temp[706] = ~window[14][2];
assign temp[707] = ~window[14][3];
assign temp[708] = ~window[14][4];
assign temp[709] = ~window[14][5];
assign temp[710] = window[14][6];
assign temp[711] = ~window[14][7];
assign temp[712] = ~window[14][8];
assign temp[736] = ~window[15][0];
assign temp[737] = window[15][1];
assign temp[738] = window[15][2];
assign temp[739] = window[15][3];
assign temp[740] = ~window[15][4];
assign temp[741] = window[15][5];
assign temp[742] = window[15][6];
assign temp[743] = window[15][7];
assign temp[744] = window[15][8];
assign temp[768] = window[16][0];
assign temp[769] = ~window[16][1];
assign temp[770] = window[16][2];
assign temp[771] = window[16][3];
assign temp[772] = window[16][4];
assign temp[773] = window[16][5];
assign temp[774] = window[16][6];
assign temp[775] = window[16][7];
assign temp[776] = window[16][8];
assign temp[800] = window[17][0];
assign temp[801] = window[17][1];
assign temp[802] = ~window[17][2];
assign temp[803] = window[17][3];
assign temp[804] = ~window[17][4];
assign temp[805] = window[17][5];
assign temp[806] = window[17][6];
assign temp[807] = window[17][7];
assign temp[808] = window[17][8];
assign temp[832] = ~window[18][0];
assign temp[833] = window[18][1];
assign temp[834] = window[18][2];
assign temp[835] = ~window[18][3];
assign temp[836] = ~window[18][4];
assign temp[837] = ~window[18][5];
assign temp[838] = window[18][6];
assign temp[839] = window[18][7];
assign temp[840] = window[18][8];
assign temp[864] = window[19][0];
assign temp[865] = window[19][1];
assign temp[866] = window[19][2];
assign temp[867] = window[19][3];
assign temp[868] = ~window[19][4];
assign temp[869] = ~window[19][5];
assign temp[870] = ~window[19][6];
assign temp[871] = ~window[19][7];
assign temp[872] = ~window[19][8];
assign temp[896] = window[20][0];
assign temp[897] = window[20][1];
assign temp[898] = ~window[20][2];
assign temp[899] = ~window[20][3];
assign temp[900] = ~window[20][4];
assign temp[901] = ~window[20][5];
assign temp[902] = window[20][6];
assign temp[903] = window[20][7];
assign temp[904] = window[20][8];
assign temp[928] = ~window[21][0];
assign temp[929] = ~window[21][1];
assign temp[930] = ~window[21][2];
assign temp[931] = window[21][3];
assign temp[932] = ~window[21][4];
assign temp[933] = window[21][5];
assign temp[934] = ~window[21][6];
assign temp[935] = ~window[21][7];
assign temp[936] = window[21][8];
assign temp[960] = ~window[22][0];
assign temp[961] = ~window[22][1];
assign temp[962] = ~window[22][2];
assign temp[963] = window[22][3];
assign temp[964] = window[22][4];
assign temp[965] = ~window[22][5];
assign temp[966] = ~window[22][6];
assign temp[967] = window[22][7];
assign temp[968] = ~window[22][8];
assign temp[992] = ~window[23][0];
assign temp[993] = ~window[23][1];
assign temp[994] = ~window[23][2];
assign temp[995] = window[23][3];
assign temp[996] = ~window[23][4];
assign temp[997] = ~window[23][5];
assign temp[998] = window[23][6];
assign temp[999] = ~window[23][7];
assign temp[1000] = window[23][8];
assign temp[1024] = window[24][0];
assign temp[1025] = window[24][1];
assign temp[1026] = ~window[24][2];
assign temp[1027] = window[24][3];
assign temp[1028] = ~window[24][4];
assign temp[1029] = ~window[24][5];
assign temp[1030] = window[24][6];
assign temp[1031] = window[24][7];
assign temp[1032] = window[24][8];
assign temp[1056] = ~window[25][0];
assign temp[1057] = window[25][1];
assign temp[1058] = window[25][2];
assign temp[1059] = ~window[25][3];
assign temp[1060] = ~window[25][4];
assign temp[1061] = ~window[25][5];
assign temp[1062] = window[25][6];
assign temp[1063] = ~window[25][7];
assign temp[1064] = window[25][8];
assign temp[1088] = ~window[26][0];
assign temp[1089] = ~window[26][1];
assign temp[1090] = ~window[26][2];
assign temp[1091] = window[26][3];
assign temp[1092] = ~window[26][4];
assign temp[1093] = window[26][5];
assign temp[1094] = ~window[26][6];
assign temp[1095] = ~window[26][7];
assign temp[1096] = ~window[26][8];
assign temp[1120] = ~window[27][0];
assign temp[1121] = ~window[27][1];
assign temp[1122] = ~window[27][2];
assign temp[1123] = window[27][3];
assign temp[1124] = window[27][4];
assign temp[1125] = ~window[27][5];
assign temp[1126] = window[27][6];
assign temp[1127] = window[27][7];
assign temp[1128] = window[27][8];
assign temp[1152] = window[28][0];
assign temp[1153] = window[28][1];
assign temp[1154] = window[28][2];
assign temp[1155] = window[28][3];
assign temp[1156] = window[28][4];
assign temp[1157] = window[28][5];
assign temp[1158] = window[28][6];
assign temp[1159] = window[28][7];
assign temp[1160] = window[28][8];
assign temp[1184] = window[29][0];
assign temp[1185] = ~window[29][1];
assign temp[1186] = ~window[29][2];
assign temp[1187] = window[29][3];
assign temp[1188] = window[29][4];
assign temp[1189] = window[29][5];
assign temp[1190] = window[29][6];
assign temp[1191] = window[29][7];
assign temp[1192] = window[29][8];
assign temp[1216] = window[30][0];
assign temp[1217] = ~window[30][1];
assign temp[1218] = ~window[30][2];
assign temp[1219] = window[30][3];
assign temp[1220] = window[30][4];
assign temp[1221] = ~window[30][5];
assign temp[1222] = window[30][6];
assign temp[1223] = ~window[30][7];
assign temp[1224] = window[30][8];
assign temp[1248] = window[31][0];
assign temp[1249] = window[31][1];
assign temp[1250] = ~window[31][2];
assign temp[1251] = window[31][3];
assign temp[1252] = window[31][4];
assign temp[1253] = ~window[31][5];
assign temp[1254] = window[31][6];
assign temp[1255] = window[31][7];
assign temp[1256] = window[31][8];
assign temp[288] = ~window[0][0];
assign temp[289] = window[0][1];
assign temp[290] = window[0][2];
assign temp[291] = window[0][3];
assign temp[292] = window[0][4];
assign temp[293] = ~window[0][5];
assign temp[294] = ~window[0][6];
assign temp[295] = ~window[0][7];
assign temp[296] = window[0][8];
assign temp[320] = ~window[1][0];
assign temp[321] = ~window[1][1];
assign temp[322] = ~window[1][2];
assign temp[323] = ~window[1][3];
assign temp[324] = ~window[1][4];
assign temp[325] = ~window[1][5];
assign temp[326] = window[1][6];
assign temp[327] = window[1][7];
assign temp[328] = window[1][8];
assign temp[352] = ~window[2][0];
assign temp[353] = window[2][1];
assign temp[354] = ~window[2][2];
assign temp[355] = ~window[2][3];
assign temp[356] = ~window[2][4];
assign temp[357] = window[2][5];
assign temp[358] = window[2][6];
assign temp[359] = window[2][7];
assign temp[360] = window[2][8];
assign temp[384] = window[3][0];
assign temp[385] = ~window[3][1];
assign temp[386] = ~window[3][2];
assign temp[387] = window[3][3];
assign temp[388] = window[3][4];
assign temp[389] = window[3][5];
assign temp[390] = window[3][6];
assign temp[391] = window[3][7];
assign temp[392] = window[3][8];
assign temp[416] = window[4][0];
assign temp[417] = ~window[4][1];
assign temp[418] = ~window[4][2];
assign temp[419] = window[4][3];
assign temp[420] = window[4][4];
assign temp[421] = window[4][5];
assign temp[422] = ~window[4][6];
assign temp[423] = ~window[4][7];
assign temp[424] = window[4][8];
assign temp[448] = ~window[5][0];
assign temp[449] = ~window[5][1];
assign temp[450] = ~window[5][2];
assign temp[451] = ~window[5][3];
assign temp[452] = ~window[5][4];
assign temp[453] = ~window[5][5];
assign temp[454] = ~window[5][6];
assign temp[455] = ~window[5][7];
assign temp[456] = ~window[5][8];
assign temp[480] = ~window[6][0];
assign temp[481] = ~window[6][1];
assign temp[482] = window[6][2];
assign temp[483] = window[6][3];
assign temp[484] = ~window[6][4];
assign temp[485] = ~window[6][5];
assign temp[486] = window[6][6];
assign temp[487] = window[6][7];
assign temp[488] = window[6][8];
assign temp[512] = window[7][0];
assign temp[513] = ~window[7][1];
assign temp[514] = ~window[7][2];
assign temp[515] = window[7][3];
assign temp[516] = window[7][4];
assign temp[517] = window[7][5];
assign temp[518] = window[7][6];
assign temp[519] = window[7][7];
assign temp[520] = ~window[7][8];
assign temp[544] = window[8][0];
assign temp[545] = ~window[8][1];
assign temp[546] = ~window[8][2];
assign temp[547] = window[8][3];
assign temp[548] = window[8][4];
assign temp[549] = window[8][5];
assign temp[550] = window[8][6];
assign temp[551] = window[8][7];
assign temp[552] = window[8][8];
assign temp[576] = ~window[9][0];
assign temp[577] = ~window[9][1];
assign temp[578] = ~window[9][2];
assign temp[579] = window[9][3];
assign temp[580] = window[9][4];
assign temp[581] = window[9][5];
assign temp[582] = window[9][6];
assign temp[583] = window[9][7];
assign temp[584] = window[9][8];
assign temp[608] = window[10][0];
assign temp[609] = ~window[10][1];
assign temp[610] = ~window[10][2];
assign temp[611] = window[10][3];
assign temp[612] = window[10][4];
assign temp[613] = window[10][5];
assign temp[614] = window[10][6];
assign temp[615] = window[10][7];
assign temp[616] = ~window[10][8];
assign temp[640] = window[11][0];
assign temp[641] = window[11][1];
assign temp[642] = window[11][2];
assign temp[643] = window[11][3];
assign temp[644] = window[11][4];
assign temp[645] = window[11][5];
assign temp[646] = ~window[11][6];
assign temp[647] = ~window[11][7];
assign temp[648] = ~window[11][8];
assign temp[672] = ~window[12][0];
assign temp[673] = window[12][1];
assign temp[674] = ~window[12][2];
assign temp[675] = ~window[12][3];
assign temp[676] = ~window[12][4];
assign temp[677] = ~window[12][5];
assign temp[678] = window[12][6];
assign temp[679] = window[12][7];
assign temp[680] = window[12][8];
assign temp[704] = ~window[13][0];
assign temp[705] = ~window[13][1];
assign temp[706] = window[13][2];
assign temp[707] = ~window[13][3];
assign temp[708] = ~window[13][4];
assign temp[709] = ~window[13][5];
assign temp[710] = ~window[13][6];
assign temp[711] = ~window[13][7];
assign temp[712] = ~window[13][8];
assign temp[736] = window[14][0];
assign temp[737] = window[14][1];
assign temp[738] = ~window[14][2];
assign temp[739] = window[14][3];
assign temp[740] = window[14][4];
assign temp[741] = window[14][5];
assign temp[742] = ~window[14][6];
assign temp[743] = ~window[14][7];
assign temp[744] = window[14][8];
assign temp[768] = window[15][0];
assign temp[769] = ~window[15][1];
assign temp[770] = window[15][2];
assign temp[771] = ~window[15][3];
assign temp[772] = window[15][4];
assign temp[773] = ~window[15][5];
assign temp[774] = window[15][6];
assign temp[775] = ~window[15][7];
assign temp[776] = ~window[15][8];
assign temp[800] = window[16][0];
assign temp[801] = ~window[16][1];
assign temp[802] = window[16][2];
assign temp[803] = window[16][3];
assign temp[804] = window[16][4];
assign temp[805] = window[16][5];
assign temp[806] = ~window[16][6];
assign temp[807] = ~window[16][7];
assign temp[808] = window[16][8];
assign temp[832] = ~window[17][0];
assign temp[833] = window[17][1];
assign temp[834] = ~window[17][2];
assign temp[835] = ~window[17][3];
assign temp[836] = ~window[17][4];
assign temp[837] = ~window[17][5];
assign temp[838] = window[17][6];
assign temp[839] = window[17][7];
assign temp[840] = window[17][8];
assign temp[864] = window[18][0];
assign temp[865] = window[18][1];
assign temp[866] = ~window[18][2];
assign temp[867] = ~window[18][3];
assign temp[868] = ~window[18][4];
assign temp[869] = ~window[18][5];
assign temp[870] = window[18][6];
assign temp[871] = window[18][7];
assign temp[872] = ~window[18][8];
assign temp[896] = ~window[19][0];
assign temp[897] = ~window[19][1];
assign temp[898] = ~window[19][2];
assign temp[899] = ~window[19][3];
assign temp[900] = ~window[19][4];
assign temp[901] = ~window[19][5];
assign temp[902] = ~window[19][6];
assign temp[903] = ~window[19][7];
assign temp[904] = ~window[19][8];
assign temp[928] = window[20][0];
assign temp[929] = ~window[20][1];
assign temp[930] = ~window[20][2];
assign temp[931] = window[20][3];
assign temp[932] = window[20][4];
assign temp[933] = window[20][5];
assign temp[934] = window[20][6];
assign temp[935] = window[20][7];
assign temp[936] = window[20][8];
assign temp[960] = window[21][0];
assign temp[961] = ~window[21][1];
assign temp[962] = ~window[21][2];
assign temp[963] = ~window[21][3];
assign temp[964] = ~window[21][4];
assign temp[965] = ~window[21][5];
assign temp[966] = ~window[21][6];
assign temp[967] = ~window[21][7];
assign temp[968] = ~window[21][8];
assign temp[992] = window[22][0];
assign temp[993] = window[22][1];
assign temp[994] = window[22][2];
assign temp[995] = ~window[22][3];
assign temp[996] = window[22][4];
assign temp[997] = ~window[22][5];
assign temp[998] = ~window[22][6];
assign temp[999] = ~window[22][7];
assign temp[1000] = ~window[22][8];
assign temp[1024] = window[23][0];
assign temp[1025] = ~window[23][1];
assign temp[1026] = ~window[23][2];
assign temp[1027] = window[23][3];
assign temp[1028] = ~window[23][4];
assign temp[1029] = ~window[23][5];
assign temp[1030] = window[23][6];
assign temp[1031] = window[23][7];
assign temp[1032] = window[23][8];
assign temp[1056] = ~window[24][0];
assign temp[1057] = window[24][1];
assign temp[1058] = window[24][2];
assign temp[1059] = ~window[24][3];
assign temp[1060] = window[24][4];
assign temp[1061] = window[24][5];
assign temp[1062] = window[24][6];
assign temp[1063] = window[24][7];
assign temp[1064] = window[24][8];
assign temp[1088] = ~window[25][0];
assign temp[1089] = ~window[25][1];
assign temp[1090] = ~window[25][2];
assign temp[1091] = ~window[25][3];
assign temp[1092] = window[25][4];
assign temp[1093] = window[25][5];
assign temp[1094] = window[25][6];
assign temp[1095] = window[25][7];
assign temp[1096] = window[25][8];
assign temp[1120] = ~window[26][0];
assign temp[1121] = ~window[26][1];
assign temp[1122] = window[26][2];
assign temp[1123] = ~window[26][3];
assign temp[1124] = ~window[26][4];
assign temp[1125] = ~window[26][5];
assign temp[1126] = ~window[26][6];
assign temp[1127] = ~window[26][7];
assign temp[1128] = ~window[26][8];
assign temp[1152] = window[27][0];
assign temp[1153] = ~window[27][1];
assign temp[1154] = ~window[27][2];
assign temp[1155] = window[27][3];
assign temp[1156] = window[27][4];
assign temp[1157] = window[27][5];
assign temp[1158] = ~window[27][6];
assign temp[1159] = ~window[27][7];
assign temp[1160] = ~window[27][8];
assign temp[1184] = window[28][0];
assign temp[1185] = window[28][1];
assign temp[1186] = window[28][2];
assign temp[1187] = window[28][3];
assign temp[1188] = ~window[28][4];
assign temp[1189] = ~window[28][5];
assign temp[1190] = window[28][6];
assign temp[1191] = window[28][7];
assign temp[1192] = ~window[28][8];
assign temp[1216] = window[29][0];
assign temp[1217] = window[29][1];
assign temp[1218] = window[29][2];
assign temp[1219] = ~window[29][3];
assign temp[1220] = window[29][4];
assign temp[1221] = window[29][5];
assign temp[1222] = ~window[29][6];
assign temp[1223] = ~window[29][7];
assign temp[1224] = ~window[29][8];
assign temp[1248] = ~window[30][0];
assign temp[1249] = ~window[30][1];
assign temp[1250] = ~window[30][2];
assign temp[1251] = ~window[30][3];
assign temp[1252] = ~window[30][4];
assign temp[1253] = ~window[30][5];
assign temp[1254] = ~window[30][6];
assign temp[1255] = ~window[30][7];
assign temp[1256] = ~window[30][8];
assign temp[1280] = ~window[31][0];
assign temp[1281] = window[31][1];
assign temp[1282] = ~window[31][2];
assign temp[1283] = window[31][3];
assign temp[1284] = window[31][4];
assign temp[1285] = window[31][5];
assign temp[1286] = window[31][6];
assign temp[1287] = window[31][7];
assign temp[1288] = window[31][8];
assign temp[320] = window[0][0];
assign temp[321] = ~window[0][1];
assign temp[322] = ~window[0][2];
assign temp[323] = ~window[0][3];
assign temp[324] = ~window[0][4];
assign temp[325] = window[0][5];
assign temp[326] = ~window[0][6];
assign temp[327] = window[0][7];
assign temp[328] = ~window[0][8];
assign temp[352] = window[1][0];
assign temp[353] = ~window[1][1];
assign temp[354] = ~window[1][2];
assign temp[355] = ~window[1][3];
assign temp[356] = ~window[1][4];
assign temp[357] = ~window[1][5];
assign temp[358] = ~window[1][6];
assign temp[359] = window[1][7];
assign temp[360] = window[1][8];
assign temp[384] = window[2][0];
assign temp[385] = ~window[2][1];
assign temp[386] = ~window[2][2];
assign temp[387] = ~window[2][3];
assign temp[388] = ~window[2][4];
assign temp[389] = window[2][5];
assign temp[390] = ~window[2][6];
assign temp[391] = ~window[2][7];
assign temp[392] = window[2][8];
assign temp[416] = window[3][0];
assign temp[417] = ~window[3][1];
assign temp[418] = ~window[3][2];
assign temp[419] = ~window[3][3];
assign temp[420] = ~window[3][4];
assign temp[421] = window[3][5];
assign temp[422] = ~window[3][6];
assign temp[423] = window[3][7];
assign temp[424] = window[3][8];
assign temp[448] = ~window[4][0];
assign temp[449] = ~window[4][1];
assign temp[450] = ~window[4][2];
assign temp[451] = ~window[4][3];
assign temp[452] = window[4][4];
assign temp[453] = ~window[4][5];
assign temp[454] = ~window[4][6];
assign temp[455] = ~window[4][7];
assign temp[456] = ~window[4][8];
assign temp[480] = window[5][0];
assign temp[481] = ~window[5][1];
assign temp[482] = ~window[5][2];
assign temp[483] = ~window[5][3];
assign temp[484] = ~window[5][4];
assign temp[485] = window[5][5];
assign temp[486] = window[5][6];
assign temp[487] = window[5][7];
assign temp[488] = ~window[5][8];
assign temp[512] = ~window[6][0];
assign temp[513] = window[6][1];
assign temp[514] = ~window[6][2];
assign temp[515] = ~window[6][3];
assign temp[516] = ~window[6][4];
assign temp[517] = ~window[6][5];
assign temp[518] = ~window[6][6];
assign temp[519] = ~window[6][7];
assign temp[520] = window[6][8];
assign temp[544] = ~window[7][0];
assign temp[545] = ~window[7][1];
assign temp[546] = ~window[7][2];
assign temp[547] = ~window[7][3];
assign temp[548] = window[7][4];
assign temp[549] = window[7][5];
assign temp[550] = window[7][6];
assign temp[551] = window[7][7];
assign temp[552] = ~window[7][8];
assign temp[576] = ~window[8][0];
assign temp[577] = ~window[8][1];
assign temp[578] = window[8][2];
assign temp[579] = ~window[8][3];
assign temp[580] = ~window[8][4];
assign temp[581] = window[8][5];
assign temp[582] = window[8][6];
assign temp[583] = window[8][7];
assign temp[584] = window[8][8];
assign temp[608] = ~window[9][0];
assign temp[609] = ~window[9][1];
assign temp[610] = ~window[9][2];
assign temp[611] = ~window[9][3];
assign temp[612] = ~window[9][4];
assign temp[613] = window[9][5];
assign temp[614] = ~window[9][6];
assign temp[615] = window[9][7];
assign temp[616] = window[9][8];
assign temp[640] = window[10][0];
assign temp[641] = ~window[10][1];
assign temp[642] = ~window[10][2];
assign temp[643] = ~window[10][3];
assign temp[644] = ~window[10][4];
assign temp[645] = ~window[10][5];
assign temp[646] = ~window[10][6];
assign temp[647] = window[10][7];
assign temp[648] = window[10][8];
assign temp[672] = window[11][0];
assign temp[673] = window[11][1];
assign temp[674] = window[11][2];
assign temp[675] = window[11][3];
assign temp[676] = ~window[11][4];
assign temp[677] = window[11][5];
assign temp[678] = window[11][6];
assign temp[679] = window[11][7];
assign temp[680] = window[11][8];
assign temp[704] = window[12][0];
assign temp[705] = window[12][1];
assign temp[706] = window[12][2];
assign temp[707] = window[12][3];
assign temp[708] = ~window[12][4];
assign temp[709] = window[12][5];
assign temp[710] = ~window[12][6];
assign temp[711] = ~window[12][7];
assign temp[712] = window[12][8];
assign temp[736] = window[13][0];
assign temp[737] = window[13][1];
assign temp[738] = window[13][2];
assign temp[739] = window[13][3];
assign temp[740] = window[13][4];
assign temp[741] = window[13][5];
assign temp[742] = ~window[13][6];
assign temp[743] = window[13][7];
assign temp[744] = window[13][8];
assign temp[768] = ~window[14][0];
assign temp[769] = ~window[14][1];
assign temp[770] = ~window[14][2];
assign temp[771] = ~window[14][3];
assign temp[772] = ~window[14][4];
assign temp[773] = ~window[14][5];
assign temp[774] = ~window[14][6];
assign temp[775] = window[14][7];
assign temp[776] = ~window[14][8];
assign temp[800] = ~window[15][0];
assign temp[801] = window[15][1];
assign temp[802] = ~window[15][2];
assign temp[803] = window[15][3];
assign temp[804] = ~window[15][4];
assign temp[805] = ~window[15][5];
assign temp[806] = ~window[15][6];
assign temp[807] = ~window[15][7];
assign temp[808] = window[15][8];
assign temp[832] = window[16][0];
assign temp[833] = window[16][1];
assign temp[834] = window[16][2];
assign temp[835] = window[16][3];
assign temp[836] = window[16][4];
assign temp[837] = window[16][5];
assign temp[838] = window[16][6];
assign temp[839] = window[16][7];
assign temp[840] = ~window[16][8];
assign temp[864] = window[17][0];
assign temp[865] = window[17][1];
assign temp[866] = ~window[17][2];
assign temp[867] = ~window[17][3];
assign temp[868] = ~window[17][4];
assign temp[869] = window[17][5];
assign temp[870] = window[17][6];
assign temp[871] = window[17][7];
assign temp[872] = window[17][8];
assign temp[896] = window[18][0];
assign temp[897] = window[18][1];
assign temp[898] = ~window[18][2];
assign temp[899] = ~window[18][3];
assign temp[900] = window[18][4];
assign temp[901] = window[18][5];
assign temp[902] = window[18][6];
assign temp[903] = ~window[18][7];
assign temp[904] = window[18][8];
assign temp[928] = window[19][0];
assign temp[929] = ~window[19][1];
assign temp[930] = ~window[19][2];
assign temp[931] = ~window[19][3];
assign temp[932] = window[19][4];
assign temp[933] = window[19][5];
assign temp[934] = ~window[19][6];
assign temp[935] = window[19][7];
assign temp[936] = ~window[19][8];
assign temp[960] = window[20][0];
assign temp[961] = ~window[20][1];
assign temp[962] = ~window[20][2];
assign temp[963] = ~window[20][3];
assign temp[964] = window[20][4];
assign temp[965] = window[20][5];
assign temp[966] = window[20][6];
assign temp[967] = window[20][7];
assign temp[968] = window[20][8];
assign temp[992] = ~window[21][0];
assign temp[993] = ~window[21][1];
assign temp[994] = ~window[21][2];
assign temp[995] = ~window[21][3];
assign temp[996] = ~window[21][4];
assign temp[997] = ~window[21][5];
assign temp[998] = ~window[21][6];
assign temp[999] = window[21][7];
assign temp[1000] = window[21][8];
assign temp[1024] = window[22][0];
assign temp[1025] = window[22][1];
assign temp[1026] = window[22][2];
assign temp[1027] = window[22][3];
assign temp[1028] = ~window[22][4];
assign temp[1029] = ~window[22][5];
assign temp[1030] = window[22][6];
assign temp[1031] = ~window[22][7];
assign temp[1032] = ~window[22][8];
assign temp[1056] = window[23][0];
assign temp[1057] = ~window[23][1];
assign temp[1058] = ~window[23][2];
assign temp[1059] = ~window[23][3];
assign temp[1060] = ~window[23][4];
assign temp[1061] = window[23][5];
assign temp[1062] = ~window[23][6];
assign temp[1063] = window[23][7];
assign temp[1064] = ~window[23][8];
assign temp[1088] = window[24][0];
assign temp[1089] = ~window[24][1];
assign temp[1090] = ~window[24][2];
assign temp[1091] = ~window[24][3];
assign temp[1092] = ~window[24][4];
assign temp[1093] = window[24][5];
assign temp[1094] = ~window[24][6];
assign temp[1095] = window[24][7];
assign temp[1096] = window[24][8];
assign temp[1120] = ~window[25][0];
assign temp[1121] = ~window[25][1];
assign temp[1122] = window[25][2];
assign temp[1123] = window[25][3];
assign temp[1124] = window[25][4];
assign temp[1125] = ~window[25][5];
assign temp[1126] = ~window[25][6];
assign temp[1127] = ~window[25][7];
assign temp[1128] = window[25][8];
assign temp[1152] = ~window[26][0];
assign temp[1153] = ~window[26][1];
assign temp[1154] = ~window[26][2];
assign temp[1155] = ~window[26][3];
assign temp[1156] = ~window[26][4];
assign temp[1157] = ~window[26][5];
assign temp[1158] = ~window[26][6];
assign temp[1159] = window[26][7];
assign temp[1160] = window[26][8];
assign temp[1184] = ~window[27][0];
assign temp[1185] = ~window[27][1];
assign temp[1186] = ~window[27][2];
assign temp[1187] = window[27][3];
assign temp[1188] = window[27][4];
assign temp[1189] = window[27][5];
assign temp[1190] = window[27][6];
assign temp[1191] = ~window[27][7];
assign temp[1192] = ~window[27][8];
assign temp[1216] = window[28][0];
assign temp[1217] = window[28][1];
assign temp[1218] = window[28][2];
assign temp[1219] = window[28][3];
assign temp[1220] = window[28][4];
assign temp[1221] = ~window[28][5];
assign temp[1222] = ~window[28][6];
assign temp[1223] = ~window[28][7];
assign temp[1224] = ~window[28][8];
assign temp[1248] = window[29][0];
assign temp[1249] = window[29][1];
assign temp[1250] = window[29][2];
assign temp[1251] = window[29][3];
assign temp[1252] = window[29][4];
assign temp[1253] = window[29][5];
assign temp[1254] = window[29][6];
assign temp[1255] = window[29][7];
assign temp[1256] = ~window[29][8];
assign temp[1280] = window[30][0];
assign temp[1281] = window[30][1];
assign temp[1282] = window[30][2];
assign temp[1283] = window[30][3];
assign temp[1284] = window[30][4];
assign temp[1285] = window[30][5];
assign temp[1286] = window[30][6];
assign temp[1287] = window[30][7];
assign temp[1288] = ~window[30][8];
assign temp[1312] = window[31][0];
assign temp[1313] = window[31][1];
assign temp[1314] = ~window[31][2];
assign temp[1315] = ~window[31][3];
assign temp[1316] = ~window[31][4];
assign temp[1317] = window[31][5];
assign temp[1318] = ~window[31][6];
assign temp[1319] = window[31][7];
assign temp[1320] = window[31][8];
assign temp[352] = window[0][0];
assign temp[353] = window[0][1];
assign temp[354] = window[0][2];
assign temp[355] = ~window[0][3];
assign temp[356] = window[0][4];
assign temp[357] = window[0][5];
assign temp[358] = window[0][6];
assign temp[359] = window[0][7];
assign temp[360] = window[0][8];
assign temp[384] = window[1][0];
assign temp[385] = window[1][1];
assign temp[386] = window[1][2];
assign temp[387] = window[1][3];
assign temp[388] = ~window[1][4];
assign temp[389] = ~window[1][5];
assign temp[390] = window[1][6];
assign temp[391] = window[1][7];
assign temp[392] = window[1][8];
assign temp[416] = window[2][0];
assign temp[417] = window[2][1];
assign temp[418] = ~window[2][2];
assign temp[419] = window[2][3];
assign temp[420] = window[2][4];
assign temp[421] = window[2][5];
assign temp[422] = window[2][6];
assign temp[423] = window[2][7];
assign temp[424] = window[2][8];
assign temp[448] = window[3][0];
assign temp[449] = window[3][1];
assign temp[450] = window[3][2];
assign temp[451] = window[3][3];
assign temp[452] = window[3][4];
assign temp[453] = window[3][5];
assign temp[454] = ~window[3][6];
assign temp[455] = ~window[3][7];
assign temp[456] = ~window[3][8];
assign temp[480] = window[4][0];
assign temp[481] = window[4][1];
assign temp[482] = window[4][2];
assign temp[483] = ~window[4][3];
assign temp[484] = ~window[4][4];
assign temp[485] = window[4][5];
assign temp[486] = ~window[4][6];
assign temp[487] = ~window[4][7];
assign temp[488] = ~window[4][8];
assign temp[512] = window[5][0];
assign temp[513] = ~window[5][1];
assign temp[514] = ~window[5][2];
assign temp[515] = ~window[5][3];
assign temp[516] = window[5][4];
assign temp[517] = window[5][5];
assign temp[518] = ~window[5][6];
assign temp[519] = ~window[5][7];
assign temp[520] = ~window[5][8];
assign temp[544] = ~window[6][0];
assign temp[545] = window[6][1];
assign temp[546] = ~window[6][2];
assign temp[547] = window[6][3];
assign temp[548] = window[6][4];
assign temp[549] = ~window[6][5];
assign temp[550] = window[6][6];
assign temp[551] = window[6][7];
assign temp[552] = window[6][8];
assign temp[576] = window[7][0];
assign temp[577] = window[7][1];
assign temp[578] = window[7][2];
assign temp[579] = ~window[7][3];
assign temp[580] = window[7][4];
assign temp[581] = window[7][5];
assign temp[582] = ~window[7][6];
assign temp[583] = ~window[7][7];
assign temp[584] = ~window[7][8];
assign temp[608] = window[8][0];
assign temp[609] = window[8][1];
assign temp[610] = window[8][2];
assign temp[611] = ~window[8][3];
assign temp[612] = ~window[8][4];
assign temp[613] = window[8][5];
assign temp[614] = ~window[8][6];
assign temp[615] = window[8][7];
assign temp[616] = window[8][8];
assign temp[640] = window[9][0];
assign temp[641] = window[9][1];
assign temp[642] = window[9][2];
assign temp[643] = ~window[9][3];
assign temp[644] = window[9][4];
assign temp[645] = ~window[9][5];
assign temp[646] = ~window[9][6];
assign temp[647] = window[9][7];
assign temp[648] = window[9][8];
assign temp[672] = window[10][0];
assign temp[673] = window[10][1];
assign temp[674] = window[10][2];
assign temp[675] = ~window[10][3];
assign temp[676] = ~window[10][4];
assign temp[677] = window[10][5];
assign temp[678] = ~window[10][6];
assign temp[679] = ~window[10][7];
assign temp[680] = ~window[10][8];
assign temp[704] = ~window[11][0];
assign temp[705] = window[11][1];
assign temp[706] = window[11][2];
assign temp[707] = ~window[11][3];
assign temp[708] = ~window[11][4];
assign temp[709] = window[11][5];
assign temp[710] = ~window[11][6];
assign temp[711] = ~window[11][7];
assign temp[712] = window[11][8];
assign temp[736] = ~window[12][0];
assign temp[737] = ~window[12][1];
assign temp[738] = window[12][2];
assign temp[739] = window[12][3];
assign temp[740] = ~window[12][4];
assign temp[741] = ~window[12][5];
assign temp[742] = window[12][6];
assign temp[743] = window[12][7];
assign temp[744] = window[12][8];
assign temp[768] = ~window[13][0];
assign temp[769] = ~window[13][1];
assign temp[770] = window[13][2];
assign temp[771] = ~window[13][3];
assign temp[772] = ~window[13][4];
assign temp[773] = window[13][5];
assign temp[774] = window[13][6];
assign temp[775] = ~window[13][7];
assign temp[776] = ~window[13][8];
assign temp[800] = window[14][0];
assign temp[801] = window[14][1];
assign temp[802] = ~window[14][2];
assign temp[803] = ~window[14][3];
assign temp[804] = ~window[14][4];
assign temp[805] = ~window[14][5];
assign temp[806] = ~window[14][6];
assign temp[807] = ~window[14][7];
assign temp[808] = ~window[14][8];
assign temp[832] = ~window[15][0];
assign temp[833] = window[15][1];
assign temp[834] = window[15][2];
assign temp[835] = window[15][3];
assign temp[836] = window[15][4];
assign temp[837] = ~window[15][5];
assign temp[838] = ~window[15][6];
assign temp[839] = window[15][7];
assign temp[840] = ~window[15][8];
assign temp[864] = window[16][0];
assign temp[865] = window[16][1];
assign temp[866] = window[16][2];
assign temp[867] = ~window[16][3];
assign temp[868] = ~window[16][4];
assign temp[869] = window[16][5];
assign temp[870] = ~window[16][6];
assign temp[871] = ~window[16][7];
assign temp[872] = ~window[16][8];
assign temp[896] = window[17][0];
assign temp[897] = window[17][1];
assign temp[898] = ~window[17][2];
assign temp[899] = ~window[17][3];
assign temp[900] = ~window[17][4];
assign temp[901] = ~window[17][5];
assign temp[902] = ~window[17][6];
assign temp[903] = window[17][7];
assign temp[904] = window[17][8];
assign temp[928] = ~window[18][0];
assign temp[929] = window[18][1];
assign temp[930] = ~window[18][2];
assign temp[931] = ~window[18][3];
assign temp[932] = ~window[18][4];
assign temp[933] = ~window[18][5];
assign temp[934] = window[18][6];
assign temp[935] = window[18][7];
assign temp[936] = window[18][8];
assign temp[960] = ~window[19][0];
assign temp[961] = ~window[19][1];
assign temp[962] = window[19][2];
assign temp[963] = ~window[19][3];
assign temp[964] = ~window[19][4];
assign temp[965] = ~window[19][5];
assign temp[966] = window[19][6];
assign temp[967] = ~window[19][7];
assign temp[968] = window[19][8];
assign temp[992] = window[20][0];
assign temp[993] = ~window[20][1];
assign temp[994] = ~window[20][2];
assign temp[995] = window[20][3];
assign temp[996] = window[20][4];
assign temp[997] = window[20][5];
assign temp[998] = ~window[20][6];
assign temp[999] = window[20][7];
assign temp[1000] = window[20][8];
assign temp[1024] = window[21][0];
assign temp[1025] = window[21][1];
assign temp[1026] = window[21][2];
assign temp[1027] = ~window[21][3];
assign temp[1028] = ~window[21][4];
assign temp[1029] = ~window[21][5];
assign temp[1030] = ~window[21][6];
assign temp[1031] = ~window[21][7];
assign temp[1032] = ~window[21][8];
assign temp[1056] = window[22][0];
assign temp[1057] = window[22][1];
assign temp[1058] = window[22][2];
assign temp[1059] = ~window[22][3];
assign temp[1060] = ~window[22][4];
assign temp[1061] = ~window[22][5];
assign temp[1062] = window[22][6];
assign temp[1063] = ~window[22][7];
assign temp[1064] = ~window[22][8];
assign temp[1088] = window[23][0];
assign temp[1089] = ~window[23][1];
assign temp[1090] = ~window[23][2];
assign temp[1091] = window[23][3];
assign temp[1092] = ~window[23][4];
assign temp[1093] = window[23][5];
assign temp[1094] = ~window[23][6];
assign temp[1095] = ~window[23][7];
assign temp[1096] = ~window[23][8];
assign temp[1120] = window[24][0];
assign temp[1121] = ~window[24][1];
assign temp[1122] = ~window[24][2];
assign temp[1123] = window[24][3];
assign temp[1124] = window[24][4];
assign temp[1125] = window[24][5];
assign temp[1126] = window[24][6];
assign temp[1127] = window[24][7];
assign temp[1128] = window[24][8];
assign temp[1152] = window[25][0];
assign temp[1153] = window[25][1];
assign temp[1154] = ~window[25][2];
assign temp[1155] = ~window[25][3];
assign temp[1156] = window[25][4];
assign temp[1157] = window[25][5];
assign temp[1158] = ~window[25][6];
assign temp[1159] = ~window[25][7];
assign temp[1160] = ~window[25][8];
assign temp[1184] = window[26][0];
assign temp[1185] = window[26][1];
assign temp[1186] = window[26][2];
assign temp[1187] = ~window[26][3];
assign temp[1188] = ~window[26][4];
assign temp[1189] = ~window[26][5];
assign temp[1190] = window[26][6];
assign temp[1191] = ~window[26][7];
assign temp[1192] = window[26][8];
assign temp[1216] = window[27][0];
assign temp[1217] = window[27][1];
assign temp[1218] = window[27][2];
assign temp[1219] = ~window[27][3];
assign temp[1220] = ~window[27][4];
assign temp[1221] = ~window[27][5];
assign temp[1222] = ~window[27][6];
assign temp[1223] = ~window[27][7];
assign temp[1224] = ~window[27][8];
assign temp[1248] = ~window[28][0];
assign temp[1249] = ~window[28][1];
assign temp[1250] = window[28][2];
assign temp[1251] = ~window[28][3];
assign temp[1252] = window[28][4];
assign temp[1253] = window[28][5];
assign temp[1254] = ~window[28][6];
assign temp[1255] = ~window[28][7];
assign temp[1256] = ~window[28][8];
assign temp[1280] = ~window[29][0];
assign temp[1281] = window[29][1];
assign temp[1282] = window[29][2];
assign temp[1283] = ~window[29][3];
assign temp[1284] = ~window[29][4];
assign temp[1285] = window[29][5];
assign temp[1286] = ~window[29][6];
assign temp[1287] = ~window[29][7];
assign temp[1288] = ~window[29][8];
assign temp[1312] = ~window[30][0];
assign temp[1313] = ~window[30][1];
assign temp[1314] = ~window[30][2];
assign temp[1315] = ~window[30][3];
assign temp[1316] = ~window[30][4];
assign temp[1317] = ~window[30][5];
assign temp[1318] = window[30][6];
assign temp[1319] = ~window[30][7];
assign temp[1320] = ~window[30][8];
assign temp[1344] = window[31][0];
assign temp[1345] = ~window[31][1];
assign temp[1346] = ~window[31][2];
assign temp[1347] = ~window[31][3];
assign temp[1348] = window[31][4];
assign temp[1349] = window[31][5];
assign temp[1350] = window[31][6];
assign temp[1351] = window[31][7];
assign temp[1352] = window[31][8];
assign temp[384] = ~window[0][0];
assign temp[385] = window[0][1];
assign temp[386] = window[0][2];
assign temp[387] = window[0][3];
assign temp[388] = window[0][4];
assign temp[389] = ~window[0][5];
assign temp[390] = window[0][6];
assign temp[391] = window[0][7];
assign temp[392] = window[0][8];
assign temp[416] = ~window[1][0];
assign temp[417] = window[1][1];
assign temp[418] = window[1][2];
assign temp[419] = window[1][3];
assign temp[420] = window[1][4];
assign temp[421] = ~window[1][5];
assign temp[422] = ~window[1][6];
assign temp[423] = ~window[1][7];
assign temp[424] = window[1][8];
assign temp[448] = window[2][0];
assign temp[449] = ~window[2][1];
assign temp[450] = window[2][2];
assign temp[451] = window[2][3];
assign temp[452] = window[2][4];
assign temp[453] = window[2][5];
assign temp[454] = window[2][6];
assign temp[455] = ~window[2][7];
assign temp[456] = window[2][8];
assign temp[480] = ~window[3][0];
assign temp[481] = window[3][1];
assign temp[482] = window[3][2];
assign temp[483] = ~window[3][3];
assign temp[484] = ~window[3][4];
assign temp[485] = window[3][5];
assign temp[486] = ~window[3][6];
assign temp[487] = ~window[3][7];
assign temp[488] = ~window[3][8];
assign temp[512] = ~window[4][0];
assign temp[513] = ~window[4][1];
assign temp[514] = window[4][2];
assign temp[515] = window[4][3];
assign temp[516] = ~window[4][4];
assign temp[517] = ~window[4][5];
assign temp[518] = window[4][6];
assign temp[519] = window[4][7];
assign temp[520] = window[4][8];
assign temp[544] = ~window[5][0];
assign temp[545] = window[5][1];
assign temp[546] = window[5][2];
assign temp[547] = window[5][3];
assign temp[548] = ~window[5][4];
assign temp[549] = window[5][5];
assign temp[550] = ~window[5][6];
assign temp[551] = ~window[5][7];
assign temp[552] = ~window[5][8];
assign temp[576] = window[6][0];
assign temp[577] = ~window[6][1];
assign temp[578] = window[6][2];
assign temp[579] = window[6][3];
assign temp[580] = window[6][4];
assign temp[581] = ~window[6][5];
assign temp[582] = ~window[6][6];
assign temp[583] = window[6][7];
assign temp[584] = window[6][8];
assign temp[608] = ~window[7][0];
assign temp[609] = ~window[7][1];
assign temp[610] = window[7][2];
assign temp[611] = ~window[7][3];
assign temp[612] = ~window[7][4];
assign temp[613] = ~window[7][5];
assign temp[614] = window[7][6];
assign temp[615] = window[7][7];
assign temp[616] = ~window[7][8];
assign temp[640] = ~window[8][0];
assign temp[641] = window[8][1];
assign temp[642] = window[8][2];
assign temp[643] = window[8][3];
assign temp[644] = window[8][4];
assign temp[645] = ~window[8][5];
assign temp[646] = ~window[8][6];
assign temp[647] = window[8][7];
assign temp[648] = window[8][8];
assign temp[672] = ~window[9][0];
assign temp[673] = window[9][1];
assign temp[674] = window[9][2];
assign temp[675] = ~window[9][3];
assign temp[676] = ~window[9][4];
assign temp[677] = window[9][5];
assign temp[678] = ~window[9][6];
assign temp[679] = ~window[9][7];
assign temp[680] = ~window[9][8];
assign temp[704] = ~window[10][0];
assign temp[705] = ~window[10][1];
assign temp[706] = ~window[10][2];
assign temp[707] = ~window[10][3];
assign temp[708] = ~window[10][4];
assign temp[709] = ~window[10][5];
assign temp[710] = ~window[10][6];
assign temp[711] = ~window[10][7];
assign temp[712] = ~window[10][8];
assign temp[736] = ~window[11][0];
assign temp[737] = ~window[11][1];
assign temp[738] = window[11][2];
assign temp[739] = window[11][3];
assign temp[740] = ~window[11][4];
assign temp[741] = ~window[11][5];
assign temp[742] = window[11][6];
assign temp[743] = ~window[11][7];
assign temp[744] = ~window[11][8];
assign temp[768] = window[12][0];
assign temp[769] = ~window[12][1];
assign temp[770] = ~window[12][2];
assign temp[771] = window[12][3];
assign temp[772] = ~window[12][4];
assign temp[773] = ~window[12][5];
assign temp[774] = ~window[12][6];
assign temp[775] = window[12][7];
assign temp[776] = window[12][8];
assign temp[800] = window[13][0];
assign temp[801] = window[13][1];
assign temp[802] = window[13][2];
assign temp[803] = ~window[13][3];
assign temp[804] = ~window[13][4];
assign temp[805] = window[13][5];
assign temp[806] = window[13][6];
assign temp[807] = ~window[13][7];
assign temp[808] = ~window[13][8];
assign temp[832] = ~window[14][0];
assign temp[833] = window[14][1];
assign temp[834] = window[14][2];
assign temp[835] = ~window[14][3];
assign temp[836] = ~window[14][4];
assign temp[837] = ~window[14][5];
assign temp[838] = window[14][6];
assign temp[839] = ~window[14][7];
assign temp[840] = ~window[14][8];
assign temp[864] = ~window[15][0];
assign temp[865] = ~window[15][1];
assign temp[866] = ~window[15][2];
assign temp[867] = window[15][3];
assign temp[868] = ~window[15][4];
assign temp[869] = ~window[15][5];
assign temp[870] = window[15][6];
assign temp[871] = window[15][7];
assign temp[872] = ~window[15][8];
assign temp[896] = ~window[16][0];
assign temp[897] = window[16][1];
assign temp[898] = window[16][2];
assign temp[899] = ~window[16][3];
assign temp[900] = ~window[16][4];
assign temp[901] = window[16][5];
assign temp[902] = window[16][6];
assign temp[903] = ~window[16][7];
assign temp[904] = ~window[16][8];
assign temp[928] = window[17][0];
assign temp[929] = window[17][1];
assign temp[930] = window[17][2];
assign temp[931] = ~window[17][3];
assign temp[932] = ~window[17][4];
assign temp[933] = window[17][5];
assign temp[934] = ~window[17][6];
assign temp[935] = ~window[17][7];
assign temp[936] = window[17][8];
assign temp[960] = ~window[18][0];
assign temp[961] = ~window[18][1];
assign temp[962] = window[18][2];
assign temp[963] = window[18][3];
assign temp[964] = window[18][4];
assign temp[965] = ~window[18][5];
assign temp[966] = ~window[18][6];
assign temp[967] = ~window[18][7];
assign temp[968] = window[18][8];
assign temp[992] = window[19][0];
assign temp[993] = window[19][1];
assign temp[994] = ~window[19][2];
assign temp[995] = window[19][3];
assign temp[996] = window[19][4];
assign temp[997] = ~window[19][5];
assign temp[998] = ~window[19][6];
assign temp[999] = window[19][7];
assign temp[1000] = window[19][8];
assign temp[1024] = window[20][0];
assign temp[1025] = window[20][1];
assign temp[1026] = window[20][2];
assign temp[1027] = ~window[20][3];
assign temp[1028] = ~window[20][4];
assign temp[1029] = window[20][5];
assign temp[1030] = ~window[20][6];
assign temp[1031] = ~window[20][7];
assign temp[1032] = ~window[20][8];
assign temp[1056] = ~window[21][0];
assign temp[1057] = window[21][1];
assign temp[1058] = window[21][2];
assign temp[1059] = window[21][3];
assign temp[1060] = ~window[21][4];
assign temp[1061] = ~window[21][5];
assign temp[1062] = window[21][6];
assign temp[1063] = window[21][7];
assign temp[1064] = window[21][8];
assign temp[1088] = ~window[22][0];
assign temp[1089] = ~window[22][1];
assign temp[1090] = ~window[22][2];
assign temp[1091] = window[22][3];
assign temp[1092] = window[22][4];
assign temp[1093] = ~window[22][5];
assign temp[1094] = window[22][6];
assign temp[1095] = window[22][7];
assign temp[1096] = window[22][8];
assign temp[1120] = window[23][0];
assign temp[1121] = window[23][1];
assign temp[1122] = window[23][2];
assign temp[1123] = ~window[23][3];
assign temp[1124] = ~window[23][4];
assign temp[1125] = window[23][5];
assign temp[1126] = ~window[23][6];
assign temp[1127] = ~window[23][7];
assign temp[1128] = ~window[23][8];
assign temp[1152] = window[24][0];
assign temp[1153] = ~window[24][1];
assign temp[1154] = window[24][2];
assign temp[1155] = window[24][3];
assign temp[1156] = window[24][4];
assign temp[1157] = window[24][5];
assign temp[1158] = ~window[24][6];
assign temp[1159] = ~window[24][7];
assign temp[1160] = window[24][8];
assign temp[1184] = window[25][0];
assign temp[1185] = window[25][1];
assign temp[1186] = window[25][2];
assign temp[1187] = ~window[25][3];
assign temp[1188] = window[25][4];
assign temp[1189] = window[25][5];
assign temp[1190] = ~window[25][6];
assign temp[1191] = ~window[25][7];
assign temp[1192] = ~window[25][8];
assign temp[1216] = ~window[26][0];
assign temp[1217] = window[26][1];
assign temp[1218] = window[26][2];
assign temp[1219] = window[26][3];
assign temp[1220] = ~window[26][4];
assign temp[1221] = ~window[26][5];
assign temp[1222] = ~window[26][6];
assign temp[1223] = window[26][7];
assign temp[1224] = window[26][8];
assign temp[1248] = ~window[27][0];
assign temp[1249] = ~window[27][1];
assign temp[1250] = window[27][2];
assign temp[1251] = ~window[27][3];
assign temp[1252] = ~window[27][4];
assign temp[1253] = ~window[27][5];
assign temp[1254] = window[27][6];
assign temp[1255] = window[27][7];
assign temp[1256] = ~window[27][8];
assign temp[1280] = ~window[28][0];
assign temp[1281] = ~window[28][1];
assign temp[1282] = window[28][2];
assign temp[1283] = ~window[28][3];
assign temp[1284] = ~window[28][4];
assign temp[1285] = ~window[28][5];
assign temp[1286] = ~window[28][6];
assign temp[1287] = ~window[28][7];
assign temp[1288] = ~window[28][8];
assign temp[1312] = ~window[29][0];
assign temp[1313] = ~window[29][1];
assign temp[1314] = window[29][2];
assign temp[1315] = ~window[29][3];
assign temp[1316] = ~window[29][4];
assign temp[1317] = window[29][5];
assign temp[1318] = window[29][6];
assign temp[1319] = window[29][7];
assign temp[1320] = window[29][8];
assign temp[1344] = window[30][0];
assign temp[1345] = ~window[30][1];
assign temp[1346] = window[30][2];
assign temp[1347] = ~window[30][3];
assign temp[1348] = ~window[30][4];
assign temp[1349] = window[30][5];
assign temp[1350] = window[30][6];
assign temp[1351] = window[30][7];
assign temp[1352] = ~window[30][8];
assign temp[1376] = window[31][0];
assign temp[1377] = ~window[31][1];
assign temp[1378] = window[31][2];
assign temp[1379] = window[31][3];
assign temp[1380] = window[31][4];
assign temp[1381] = window[31][5];
assign temp[1382] = window[31][6];
assign temp[1383] = ~window[31][7];
assign temp[1384] = window[31][8];
assign temp[416] = ~window[0][0];
assign temp[417] = ~window[0][1];
assign temp[418] = window[0][2];
assign temp[419] = window[0][3];
assign temp[420] = window[0][4];
assign temp[421] = ~window[0][5];
assign temp[422] = ~window[0][6];
assign temp[423] = ~window[0][7];
assign temp[424] = ~window[0][8];
assign temp[448] = window[1][0];
assign temp[449] = window[1][1];
assign temp[450] = window[1][2];
assign temp[451] = ~window[1][3];
assign temp[452] = ~window[1][4];
assign temp[453] = ~window[1][5];
assign temp[454] = ~window[1][6];
assign temp[455] = ~window[1][7];
assign temp[456] = ~window[1][8];
assign temp[480] = window[2][0];
assign temp[481] = window[2][1];
assign temp[482] = window[2][2];
assign temp[483] = window[2][3];
assign temp[484] = window[2][4];
assign temp[485] = window[2][5];
assign temp[486] = window[2][6];
assign temp[487] = window[2][7];
assign temp[488] = ~window[2][8];
assign temp[512] = window[3][0];
assign temp[513] = window[3][1];
assign temp[514] = window[3][2];
assign temp[515] = ~window[3][3];
assign temp[516] = ~window[3][4];
assign temp[517] = ~window[3][5];
assign temp[518] = ~window[3][6];
assign temp[519] = ~window[3][7];
assign temp[520] = window[3][8];
assign temp[544] = ~window[4][0];
assign temp[545] = window[4][1];
assign temp[546] = ~window[4][2];
assign temp[547] = ~window[4][3];
assign temp[548] = ~window[4][4];
assign temp[549] = ~window[4][5];
assign temp[550] = window[4][6];
assign temp[551] = window[4][7];
assign temp[552] = window[4][8];
assign temp[576] = ~window[5][0];
assign temp[577] = window[5][1];
assign temp[578] = ~window[5][2];
assign temp[579] = ~window[5][3];
assign temp[580] = ~window[5][4];
assign temp[581] = ~window[5][5];
assign temp[582] = ~window[5][6];
assign temp[583] = ~window[5][7];
assign temp[584] = window[5][8];
assign temp[608] = ~window[6][0];
assign temp[609] = ~window[6][1];
assign temp[610] = ~window[6][2];
assign temp[611] = window[6][3];
assign temp[612] = window[6][4];
assign temp[613] = window[6][5];
assign temp[614] = ~window[6][6];
assign temp[615] = ~window[6][7];
assign temp[616] = ~window[6][8];
assign temp[640] = window[7][0];
assign temp[641] = ~window[7][1];
assign temp[642] = ~window[7][2];
assign temp[643] = ~window[7][3];
assign temp[644] = ~window[7][4];
assign temp[645] = ~window[7][5];
assign temp[646] = ~window[7][6];
assign temp[647] = window[7][7];
assign temp[648] = window[7][8];
assign temp[672] = ~window[8][0];
assign temp[673] = ~window[8][1];
assign temp[674] = ~window[8][2];
assign temp[675] = window[8][3];
assign temp[676] = window[8][4];
assign temp[677] = ~window[8][5];
assign temp[678] = window[8][6];
assign temp[679] = window[8][7];
assign temp[680] = window[8][8];
assign temp[704] = window[9][0];
assign temp[705] = window[9][1];
assign temp[706] = window[9][2];
assign temp[707] = ~window[9][3];
assign temp[708] = ~window[9][4];
assign temp[709] = ~window[9][5];
assign temp[710] = ~window[9][6];
assign temp[711] = window[9][7];
assign temp[712] = ~window[9][8];
assign temp[736] = window[10][0];
assign temp[737] = ~window[10][1];
assign temp[738] = window[10][2];
assign temp[739] = ~window[10][3];
assign temp[740] = ~window[10][4];
assign temp[741] = ~window[10][5];
assign temp[742] = ~window[10][6];
assign temp[743] = ~window[10][7];
assign temp[744] = ~window[10][8];
assign temp[768] = window[11][0];
assign temp[769] = ~window[11][1];
assign temp[770] = ~window[11][2];
assign temp[771] = window[11][3];
assign temp[772] = window[11][4];
assign temp[773] = window[11][5];
assign temp[774] = window[11][6];
assign temp[775] = window[11][7];
assign temp[776] = ~window[11][8];
assign temp[800] = ~window[12][0];
assign temp[801] = ~window[12][1];
assign temp[802] = ~window[12][2];
assign temp[803] = window[12][3];
assign temp[804] = window[12][4];
assign temp[805] = window[12][5];
assign temp[806] = window[12][6];
assign temp[807] = window[12][7];
assign temp[808] = ~window[12][8];
assign temp[832] = ~window[13][0];
assign temp[833] = ~window[13][1];
assign temp[834] = window[13][2];
assign temp[835] = ~window[13][3];
assign temp[836] = window[13][4];
assign temp[837] = window[13][5];
assign temp[838] = window[13][6];
assign temp[839] = window[13][7];
assign temp[840] = ~window[13][8];
assign temp[864] = ~window[14][0];
assign temp[865] = ~window[14][1];
assign temp[866] = ~window[14][2];
assign temp[867] = ~window[14][3];
assign temp[868] = window[14][4];
assign temp[869] = ~window[14][5];
assign temp[870] = window[14][6];
assign temp[871] = window[14][7];
assign temp[872] = window[14][8];
assign temp[896] = window[15][0];
assign temp[897] = ~window[15][1];
assign temp[898] = ~window[15][2];
assign temp[899] = ~window[15][3];
assign temp[900] = ~window[15][4];
assign temp[901] = ~window[15][5];
assign temp[902] = ~window[15][6];
assign temp[903] = window[15][7];
assign temp[904] = ~window[15][8];
assign temp[928] = ~window[16][0];
assign temp[929] = ~window[16][1];
assign temp[930] = ~window[16][2];
assign temp[931] = ~window[16][3];
assign temp[932] = ~window[16][4];
assign temp[933] = ~window[16][5];
assign temp[934] = window[16][6];
assign temp[935] = window[16][7];
assign temp[936] = window[16][8];
assign temp[960] = window[17][0];
assign temp[961] = window[17][1];
assign temp[962] = window[17][2];
assign temp[963] = ~window[17][3];
assign temp[964] = ~window[17][4];
assign temp[965] = ~window[17][5];
assign temp[966] = ~window[17][6];
assign temp[967] = ~window[17][7];
assign temp[968] = ~window[17][8];
assign temp[992] = ~window[18][0];
assign temp[993] = window[18][1];
assign temp[994] = window[18][2];
assign temp[995] = ~window[18][3];
assign temp[996] = ~window[18][4];
assign temp[997] = ~window[18][5];
assign temp[998] = ~window[18][6];
assign temp[999] = ~window[18][7];
assign temp[1000] = window[18][8];
assign temp[1024] = ~window[19][0];
assign temp[1025] = window[19][1];
assign temp[1026] = window[19][2];
assign temp[1027] = ~window[19][3];
assign temp[1028] = ~window[19][4];
assign temp[1029] = window[19][5];
assign temp[1030] = window[19][6];
assign temp[1031] = ~window[19][7];
assign temp[1032] = ~window[19][8];
assign temp[1056] = ~window[20][0];
assign temp[1057] = window[20][1];
assign temp[1058] = window[20][2];
assign temp[1059] = ~window[20][3];
assign temp[1060] = ~window[20][4];
assign temp[1061] = ~window[20][5];
assign temp[1062] = ~window[20][6];
assign temp[1063] = window[20][7];
assign temp[1064] = ~window[20][8];
assign temp[1088] = ~window[21][0];
assign temp[1089] = window[21][1];
assign temp[1090] = ~window[21][2];
assign temp[1091] = ~window[21][3];
assign temp[1092] = ~window[21][4];
assign temp[1093] = ~window[21][5];
assign temp[1094] = ~window[21][6];
assign temp[1095] = ~window[21][7];
assign temp[1096] = ~window[21][8];
assign temp[1120] = ~window[22][0];
assign temp[1121] = window[22][1];
assign temp[1122] = ~window[22][2];
assign temp[1123] = window[22][3];
assign temp[1124] = ~window[22][4];
assign temp[1125] = window[22][5];
assign temp[1126] = window[22][6];
assign temp[1127] = window[22][7];
assign temp[1128] = window[22][8];
assign temp[1152] = window[23][0];
assign temp[1153] = window[23][1];
assign temp[1154] = ~window[23][2];
assign temp[1155] = ~window[23][3];
assign temp[1156] = ~window[23][4];
assign temp[1157] = ~window[23][5];
assign temp[1158] = ~window[23][6];
assign temp[1159] = window[23][7];
assign temp[1160] = ~window[23][8];
assign temp[1184] = ~window[24][0];
assign temp[1185] = ~window[24][1];
assign temp[1186] = window[24][2];
assign temp[1187] = window[24][3];
assign temp[1188] = window[24][4];
assign temp[1189] = ~window[24][5];
assign temp[1190] = ~window[24][6];
assign temp[1191] = ~window[24][7];
assign temp[1192] = ~window[24][8];
assign temp[1216] = ~window[25][0];
assign temp[1217] = window[25][1];
assign temp[1218] = ~window[25][2];
assign temp[1219] = ~window[25][3];
assign temp[1220] = ~window[25][4];
assign temp[1221] = ~window[25][5];
assign temp[1222] = window[25][6];
assign temp[1223] = window[25][7];
assign temp[1224] = ~window[25][8];
assign temp[1248] = window[26][0];
assign temp[1249] = ~window[26][1];
assign temp[1250] = ~window[26][2];
assign temp[1251] = ~window[26][3];
assign temp[1252] = window[26][4];
assign temp[1253] = window[26][5];
assign temp[1254] = ~window[26][6];
assign temp[1255] = ~window[26][7];
assign temp[1256] = ~window[26][8];
assign temp[1280] = ~window[27][0];
assign temp[1281] = ~window[27][1];
assign temp[1282] = ~window[27][2];
assign temp[1283] = ~window[27][3];
assign temp[1284] = ~window[27][4];
assign temp[1285] = ~window[27][5];
assign temp[1286] = ~window[27][6];
assign temp[1287] = window[27][7];
assign temp[1288] = window[27][8];
assign temp[1312] = ~window[28][0];
assign temp[1313] = ~window[28][1];
assign temp[1314] = ~window[28][2];
assign temp[1315] = window[28][3];
assign temp[1316] = window[28][4];
assign temp[1317] = window[28][5];
assign temp[1318] = window[28][6];
assign temp[1319] = window[28][7];
assign temp[1320] = window[28][8];
assign temp[1344] = window[29][0];
assign temp[1345] = ~window[29][1];
assign temp[1346] = ~window[29][2];
assign temp[1347] = window[29][3];
assign temp[1348] = window[29][4];
assign temp[1349] = window[29][5];
assign temp[1350] = window[29][6];
assign temp[1351] = window[29][7];
assign temp[1352] = window[29][8];
assign temp[1376] = ~window[30][0];
assign temp[1377] = ~window[30][1];
assign temp[1378] = window[30][2];
assign temp[1379] = window[30][3];
assign temp[1380] = ~window[30][4];
assign temp[1381] = ~window[30][5];
assign temp[1382] = window[30][6];
assign temp[1383] = window[30][7];
assign temp[1384] = ~window[30][8];
assign temp[1408] = window[31][0];
assign temp[1409] = window[31][1];
assign temp[1410] = window[31][2];
assign temp[1411] = window[31][3];
assign temp[1412] = window[31][4];
assign temp[1413] = window[31][5];
assign temp[1414] = window[31][6];
assign temp[1415] = window[31][7];
assign temp[1416] = window[31][8];
assign temp[448] = window[0][0];
assign temp[449] = ~window[0][1];
assign temp[450] = ~window[0][2];
assign temp[451] = ~window[0][3];
assign temp[452] = ~window[0][4];
assign temp[453] = ~window[0][5];
assign temp[454] = window[0][6];
assign temp[455] = window[0][7];
assign temp[456] = window[0][8];
assign temp[480] = window[1][0];
assign temp[481] = window[1][1];
assign temp[482] = ~window[1][2];
assign temp[483] = window[1][3];
assign temp[484] = window[1][4];
assign temp[485] = ~window[1][5];
assign temp[486] = window[1][6];
assign temp[487] = window[1][7];
assign temp[488] = window[1][8];
assign temp[512] = ~window[2][0];
assign temp[513] = ~window[2][1];
assign temp[514] = ~window[2][2];
assign temp[515] = window[2][3];
assign temp[516] = ~window[2][4];
assign temp[517] = ~window[2][5];
assign temp[518] = ~window[2][6];
assign temp[519] = ~window[2][7];
assign temp[520] = window[2][8];
assign temp[544] = window[3][0];
assign temp[545] = window[3][1];
assign temp[546] = ~window[3][2];
assign temp[547] = window[3][3];
assign temp[548] = window[3][4];
assign temp[549] = window[3][5];
assign temp[550] = ~window[3][6];
assign temp[551] = window[3][7];
assign temp[552] = window[3][8];
assign temp[576] = window[4][0];
assign temp[577] = ~window[4][1];
assign temp[578] = ~window[4][2];
assign temp[579] = ~window[4][3];
assign temp[580] = ~window[4][4];
assign temp[581] = window[4][5];
assign temp[582] = window[4][6];
assign temp[583] = window[4][7];
assign temp[584] = window[4][8];
assign temp[608] = window[5][0];
assign temp[609] = ~window[5][1];
assign temp[610] = ~window[5][2];
assign temp[611] = ~window[5][3];
assign temp[612] = ~window[5][4];
assign temp[613] = window[5][5];
assign temp[614] = ~window[5][6];
assign temp[615] = window[5][7];
assign temp[616] = window[5][8];
assign temp[640] = ~window[6][0];
assign temp[641] = ~window[6][1];
assign temp[642] = ~window[6][2];
assign temp[643] = ~window[6][3];
assign temp[644] = window[6][4];
assign temp[645] = ~window[6][5];
assign temp[646] = ~window[6][6];
assign temp[647] = ~window[6][7];
assign temp[648] = ~window[6][8];
assign temp[672] = window[7][0];
assign temp[673] = window[7][1];
assign temp[674] = ~window[7][2];
assign temp[675] = ~window[7][3];
assign temp[676] = window[7][4];
assign temp[677] = window[7][5];
assign temp[678] = ~window[7][6];
assign temp[679] = window[7][7];
assign temp[680] = window[7][8];
assign temp[704] = ~window[8][0];
assign temp[705] = ~window[8][1];
assign temp[706] = ~window[8][2];
assign temp[707] = window[8][3];
assign temp[708] = window[8][4];
assign temp[709] = window[8][5];
assign temp[710] = window[8][6];
assign temp[711] = window[8][7];
assign temp[712] = window[8][8];
assign temp[736] = window[9][0];
assign temp[737] = window[9][1];
assign temp[738] = window[9][2];
assign temp[739] = window[9][3];
assign temp[740] = window[9][4];
assign temp[741] = window[9][5];
assign temp[742] = window[9][6];
assign temp[743] = window[9][7];
assign temp[744] = window[9][8];
assign temp[768] = window[10][0];
assign temp[769] = window[10][1];
assign temp[770] = ~window[10][2];
assign temp[771] = window[10][3];
assign temp[772] = ~window[10][4];
assign temp[773] = window[10][5];
assign temp[774] = ~window[10][6];
assign temp[775] = window[10][7];
assign temp[776] = window[10][8];
assign temp[800] = window[11][0];
assign temp[801] = window[11][1];
assign temp[802] = window[11][2];
assign temp[803] = window[11][3];
assign temp[804] = ~window[11][4];
assign temp[805] = ~window[11][5];
assign temp[806] = ~window[11][6];
assign temp[807] = ~window[11][7];
assign temp[808] = ~window[11][8];
assign temp[832] = ~window[12][0];
assign temp[833] = ~window[12][1];
assign temp[834] = window[12][2];
assign temp[835] = window[12][3];
assign temp[836] = ~window[12][4];
assign temp[837] = window[12][5];
assign temp[838] = window[12][6];
assign temp[839] = ~window[12][7];
assign temp[840] = ~window[12][8];
assign temp[864] = ~window[13][0];
assign temp[865] = ~window[13][1];
assign temp[866] = window[13][2];
assign temp[867] = window[13][3];
assign temp[868] = window[13][4];
assign temp[869] = window[13][5];
assign temp[870] = window[13][6];
assign temp[871] = window[13][7];
assign temp[872] = window[13][8];
assign temp[896] = window[14][0];
assign temp[897] = window[14][1];
assign temp[898] = window[14][2];
assign temp[899] = ~window[14][3];
assign temp[900] = window[14][4];
assign temp[901] = window[14][5];
assign temp[902] = window[14][6];
assign temp[903] = window[14][7];
assign temp[904] = window[14][8];
assign temp[928] = ~window[15][0];
assign temp[929] = window[15][1];
assign temp[930] = window[15][2];
assign temp[931] = window[15][3];
assign temp[932] = ~window[15][4];
assign temp[933] = ~window[15][5];
assign temp[934] = ~window[15][6];
assign temp[935] = ~window[15][7];
assign temp[936] = window[15][8];
assign temp[960] = ~window[16][0];
assign temp[961] = ~window[16][1];
assign temp[962] = window[16][2];
assign temp[963] = ~window[16][3];
assign temp[964] = window[16][4];
assign temp[965] = window[16][5];
assign temp[966] = window[16][6];
assign temp[967] = window[16][7];
assign temp[968] = window[16][8];
assign temp[992] = window[17][0];
assign temp[993] = window[17][1];
assign temp[994] = ~window[17][2];
assign temp[995] = window[17][3];
assign temp[996] = ~window[17][4];
assign temp[997] = ~window[17][5];
assign temp[998] = ~window[17][6];
assign temp[999] = window[17][7];
assign temp[1000] = window[17][8];
assign temp[1024] = ~window[18][0];
assign temp[1025] = window[18][1];
assign temp[1026] = ~window[18][2];
assign temp[1027] = window[18][3];
assign temp[1028] = window[18][4];
assign temp[1029] = window[18][5];
assign temp[1030] = window[18][6];
assign temp[1031] = window[18][7];
assign temp[1032] = window[18][8];
assign temp[1056] = ~window[19][0];
assign temp[1057] = window[19][1];
assign temp[1058] = window[19][2];
assign temp[1059] = window[19][3];
assign temp[1060] = window[19][4];
assign temp[1061] = ~window[19][5];
assign temp[1062] = ~window[19][6];
assign temp[1063] = ~window[19][7];
assign temp[1064] = window[19][8];
assign temp[1088] = window[20][0];
assign temp[1089] = window[20][1];
assign temp[1090] = window[20][2];
assign temp[1091] = window[20][3];
assign temp[1092] = window[20][4];
assign temp[1093] = window[20][5];
assign temp[1094] = ~window[20][6];
assign temp[1095] = window[20][7];
assign temp[1096] = window[20][8];
assign temp[1120] = window[21][0];
assign temp[1121] = window[21][1];
assign temp[1122] = window[21][2];
assign temp[1123] = ~window[21][3];
assign temp[1124] = window[21][4];
assign temp[1125] = ~window[21][5];
assign temp[1126] = window[21][6];
assign temp[1127] = window[21][7];
assign temp[1128] = window[21][8];
assign temp[1152] = ~window[22][0];
assign temp[1153] = ~window[22][1];
assign temp[1154] = window[22][2];
assign temp[1155] = ~window[22][3];
assign temp[1156] = ~window[22][4];
assign temp[1157] = ~window[22][5];
assign temp[1158] = ~window[22][6];
assign temp[1159] = ~window[22][7];
assign temp[1160] = ~window[22][8];
assign temp[1184] = window[23][0];
assign temp[1185] = window[23][1];
assign temp[1186] = ~window[23][2];
assign temp[1187] = window[23][3];
assign temp[1188] = ~window[23][4];
assign temp[1189] = ~window[23][5];
assign temp[1190] = ~window[23][6];
assign temp[1191] = window[23][7];
assign temp[1192] = window[23][8];
assign temp[1216] = window[24][0];
assign temp[1217] = ~window[24][1];
assign temp[1218] = ~window[24][2];
assign temp[1219] = window[24][3];
assign temp[1220] = ~window[24][4];
assign temp[1221] = ~window[24][5];
assign temp[1222] = window[24][6];
assign temp[1223] = ~window[24][7];
assign temp[1224] = window[24][8];
assign temp[1248] = window[25][0];
assign temp[1249] = ~window[25][1];
assign temp[1250] = window[25][2];
assign temp[1251] = ~window[25][3];
assign temp[1252] = ~window[25][4];
assign temp[1253] = window[25][5];
assign temp[1254] = window[25][6];
assign temp[1255] = window[25][7];
assign temp[1256] = window[25][8];
assign temp[1280] = ~window[26][0];
assign temp[1281] = ~window[26][1];
assign temp[1282] = ~window[26][2];
assign temp[1283] = ~window[26][3];
assign temp[1284] = ~window[26][4];
assign temp[1285] = ~window[26][5];
assign temp[1286] = ~window[26][6];
assign temp[1287] = ~window[26][7];
assign temp[1288] = ~window[26][8];
assign temp[1312] = window[27][0];
assign temp[1313] = window[27][1];
assign temp[1314] = window[27][2];
assign temp[1315] = ~window[27][3];
assign temp[1316] = ~window[27][4];
assign temp[1317] = window[27][5];
assign temp[1318] = window[27][6];
assign temp[1319] = window[27][7];
assign temp[1320] = window[27][8];
assign temp[1344] = ~window[28][0];
assign temp[1345] = ~window[28][1];
assign temp[1346] = window[28][2];
assign temp[1347] = window[28][3];
assign temp[1348] = window[28][4];
assign temp[1349] = window[28][5];
assign temp[1350] = window[28][6];
assign temp[1351] = window[28][7];
assign temp[1352] = window[28][8];
assign temp[1376] = window[29][0];
assign temp[1377] = ~window[29][1];
assign temp[1378] = window[29][2];
assign temp[1379] = ~window[29][3];
assign temp[1380] = window[29][4];
assign temp[1381] = window[29][5];
assign temp[1382] = window[29][6];
assign temp[1383] = window[29][7];
assign temp[1384] = window[29][8];
assign temp[1408] = ~window[30][0];
assign temp[1409] = ~window[30][1];
assign temp[1410] = ~window[30][2];
assign temp[1411] = ~window[30][3];
assign temp[1412] = ~window[30][4];
assign temp[1413] = window[30][5];
assign temp[1414] = window[30][6];
assign temp[1415] = window[30][7];
assign temp[1416] = window[30][8];
assign temp[1440] = ~window[31][0];
assign temp[1441] = ~window[31][1];
assign temp[1442] = window[31][2];
assign temp[1443] = window[31][3];
assign temp[1444] = ~window[31][4];
assign temp[1445] = ~window[31][5];
assign temp[1446] = ~window[31][6];
assign temp[1447] = window[31][7];
assign temp[1448] = window[31][8];
assign temp[480] = ~window[0][0];
assign temp[481] = ~window[0][1];
assign temp[482] = ~window[0][2];
assign temp[483] = ~window[0][3];
assign temp[484] = window[0][4];
assign temp[485] = ~window[0][5];
assign temp[486] = window[0][6];
assign temp[487] = window[0][7];
assign temp[488] = ~window[0][8];
assign temp[512] = window[1][0];
assign temp[513] = window[1][1];
assign temp[514] = window[1][2];
assign temp[515] = ~window[1][3];
assign temp[516] = window[1][4];
assign temp[517] = ~window[1][5];
assign temp[518] = window[1][6];
assign temp[519] = window[1][7];
assign temp[520] = window[1][8];
assign temp[544] = ~window[2][0];
assign temp[545] = ~window[2][1];
assign temp[546] = ~window[2][2];
assign temp[547] = window[2][3];
assign temp[548] = ~window[2][4];
assign temp[549] = ~window[2][5];
assign temp[550] = ~window[2][6];
assign temp[551] = ~window[2][7];
assign temp[552] = ~window[2][8];
assign temp[576] = window[3][0];
assign temp[577] = ~window[3][1];
assign temp[578] = ~window[3][2];
assign temp[579] = window[3][3];
assign temp[580] = ~window[3][4];
assign temp[581] = ~window[3][5];
assign temp[582] = window[3][6];
assign temp[583] = ~window[3][7];
assign temp[584] = window[3][8];
assign temp[608] = window[4][0];
assign temp[609] = ~window[4][1];
assign temp[610] = ~window[4][2];
assign temp[611] = ~window[4][3];
assign temp[612] = window[4][4];
assign temp[613] = window[4][5];
assign temp[614] = window[4][6];
assign temp[615] = window[4][7];
assign temp[616] = window[4][8];
assign temp[640] = window[5][0];
assign temp[641] = ~window[5][1];
assign temp[642] = window[5][2];
assign temp[643] = window[5][3];
assign temp[644] = window[5][4];
assign temp[645] = window[5][5];
assign temp[646] = window[5][6];
assign temp[647] = window[5][7];
assign temp[648] = ~window[5][8];
assign temp[672] = ~window[6][0];
assign temp[673] = ~window[6][1];
assign temp[674] = window[6][2];
assign temp[675] = ~window[6][3];
assign temp[676] = window[6][4];
assign temp[677] = ~window[6][5];
assign temp[678] = window[6][6];
assign temp[679] = window[6][7];
assign temp[680] = ~window[6][8];
assign temp[704] = window[7][0];
assign temp[705] = window[7][1];
assign temp[706] = ~window[7][2];
assign temp[707] = window[7][3];
assign temp[708] = window[7][4];
assign temp[709] = ~window[7][5];
assign temp[710] = ~window[7][6];
assign temp[711] = window[7][7];
assign temp[712] = window[7][8];
assign temp[736] = ~window[8][0];
assign temp[737] = ~window[8][1];
assign temp[738] = ~window[8][2];
assign temp[739] = ~window[8][3];
assign temp[740] = ~window[8][4];
assign temp[741] = ~window[8][5];
assign temp[742] = ~window[8][6];
assign temp[743] = window[8][7];
assign temp[744] = ~window[8][8];
assign temp[768] = window[9][0];
assign temp[769] = window[9][1];
assign temp[770] = ~window[9][2];
assign temp[771] = window[9][3];
assign temp[772] = window[9][4];
assign temp[773] = ~window[9][5];
assign temp[774] = ~window[9][6];
assign temp[775] = window[9][7];
assign temp[776] = ~window[9][8];
assign temp[800] = window[10][0];
assign temp[801] = window[10][1];
assign temp[802] = ~window[10][2];
assign temp[803] = window[10][3];
assign temp[804] = window[10][4];
assign temp[805] = ~window[10][5];
assign temp[806] = window[10][6];
assign temp[807] = window[10][7];
assign temp[808] = window[10][8];
assign temp[832] = window[11][0];
assign temp[833] = window[11][1];
assign temp[834] = ~window[11][2];
assign temp[835] = ~window[11][3];
assign temp[836] = ~window[11][4];
assign temp[837] = ~window[11][5];
assign temp[838] = ~window[11][6];
assign temp[839] = ~window[11][7];
assign temp[840] = ~window[11][8];
assign temp[864] = ~window[12][0];
assign temp[865] = ~window[12][1];
assign temp[866] = window[12][2];
assign temp[867] = ~window[12][3];
assign temp[868] = ~window[12][4];
assign temp[869] = ~window[12][5];
assign temp[870] = ~window[12][6];
assign temp[871] = ~window[12][7];
assign temp[872] = window[12][8];
assign temp[896] = window[13][0];
assign temp[897] = ~window[13][1];
assign temp[898] = window[13][2];
assign temp[899] = window[13][3];
assign temp[900] = ~window[13][4];
assign temp[901] = window[13][5];
assign temp[902] = window[13][6];
assign temp[903] = ~window[13][7];
assign temp[904] = window[13][8];
assign temp[928] = ~window[14][0];
assign temp[929] = ~window[14][1];
assign temp[930] = ~window[14][2];
assign temp[931] = window[14][3];
assign temp[932] = ~window[14][4];
assign temp[933] = ~window[14][5];
assign temp[934] = window[14][6];
assign temp[935] = ~window[14][7];
assign temp[936] = ~window[14][8];
assign temp[960] = ~window[15][0];
assign temp[961] = window[15][1];
assign temp[962] = ~window[15][2];
assign temp[963] = ~window[15][3];
assign temp[964] = window[15][4];
assign temp[965] = window[15][5];
assign temp[966] = ~window[15][6];
assign temp[967] = window[15][7];
assign temp[968] = window[15][8];
assign temp[992] = window[16][0];
assign temp[993] = ~window[16][1];
assign temp[994] = ~window[16][2];
assign temp[995] = window[16][3];
assign temp[996] = window[16][4];
assign temp[997] = ~window[16][5];
assign temp[998] = window[16][6];
assign temp[999] = ~window[16][7];
assign temp[1000] = window[16][8];
assign temp[1024] = window[17][0];
assign temp[1025] = window[17][1];
assign temp[1026] = ~window[17][2];
assign temp[1027] = ~window[17][3];
assign temp[1028] = window[17][4];
assign temp[1029] = ~window[17][5];
assign temp[1030] = window[17][6];
assign temp[1031] = window[17][7];
assign temp[1032] = ~window[17][8];
assign temp[1056] = ~window[18][0];
assign temp[1057] = ~window[18][1];
assign temp[1058] = window[18][2];
assign temp[1059] = window[18][3];
assign temp[1060] = ~window[18][4];
assign temp[1061] = window[18][5];
assign temp[1062] = window[18][6];
assign temp[1063] = ~window[18][7];
assign temp[1064] = ~window[18][8];
assign temp[1088] = window[19][0];
assign temp[1089] = window[19][1];
assign temp[1090] = window[19][2];
assign temp[1091] = ~window[19][3];
assign temp[1092] = ~window[19][4];
assign temp[1093] = window[19][5];
assign temp[1094] = window[19][6];
assign temp[1095] = ~window[19][7];
assign temp[1096] = window[19][8];
assign temp[1120] = window[20][0];
assign temp[1121] = window[20][1];
assign temp[1122] = ~window[20][2];
assign temp[1123] = window[20][3];
assign temp[1124] = window[20][4];
assign temp[1125] = ~window[20][5];
assign temp[1126] = window[20][6];
assign temp[1127] = ~window[20][7];
assign temp[1128] = ~window[20][8];
assign temp[1152] = window[21][0];
assign temp[1153] = window[21][1];
assign temp[1154] = window[21][2];
assign temp[1155] = window[21][3];
assign temp[1156] = window[21][4];
assign temp[1157] = window[21][5];
assign temp[1158] = window[21][6];
assign temp[1159] = window[21][7];
assign temp[1160] = window[21][8];
assign temp[1184] = ~window[22][0];
assign temp[1185] = ~window[22][1];
assign temp[1186] = window[22][2];
assign temp[1187] = ~window[22][3];
assign temp[1188] = window[22][4];
assign temp[1189] = window[22][5];
assign temp[1190] = ~window[22][6];
assign temp[1191] = ~window[22][7];
assign temp[1192] = window[22][8];
assign temp[1216] = window[23][0];
assign temp[1217] = ~window[23][1];
assign temp[1218] = window[23][2];
assign temp[1219] = window[23][3];
assign temp[1220] = ~window[23][4];
assign temp[1221] = window[23][5];
assign temp[1222] = window[23][6];
assign temp[1223] = window[23][7];
assign temp[1224] = window[23][8];
assign temp[1248] = ~window[24][0];
assign temp[1249] = ~window[24][1];
assign temp[1250] = window[24][2];
assign temp[1251] = window[24][3];
assign temp[1252] = ~window[24][4];
assign temp[1253] = ~window[24][5];
assign temp[1254] = ~window[24][6];
assign temp[1255] = ~window[24][7];
assign temp[1256] = ~window[24][8];
assign temp[1280] = window[25][0];
assign temp[1281] = ~window[25][1];
assign temp[1282] = window[25][2];
assign temp[1283] = window[25][3];
assign temp[1284] = ~window[25][4];
assign temp[1285] = ~window[25][5];
assign temp[1286] = ~window[25][6];
assign temp[1287] = ~window[25][7];
assign temp[1288] = ~window[25][8];
assign temp[1312] = window[26][0];
assign temp[1313] = window[26][1];
assign temp[1314] = window[26][2];
assign temp[1315] = window[26][3];
assign temp[1316] = window[26][4];
assign temp[1317] = window[26][5];
assign temp[1318] = ~window[26][6];
assign temp[1319] = ~window[26][7];
assign temp[1320] = window[26][8];
assign temp[1344] = window[27][0];
assign temp[1345] = ~window[27][1];
assign temp[1346] = ~window[27][2];
assign temp[1347] = ~window[27][3];
assign temp[1348] = window[27][4];
assign temp[1349] = window[27][5];
assign temp[1350] = ~window[27][6];
assign temp[1351] = window[27][7];
assign temp[1352] = ~window[27][8];
assign temp[1376] = window[28][0];
assign temp[1377] = window[28][1];
assign temp[1378] = window[28][2];
assign temp[1379] = window[28][3];
assign temp[1380] = window[28][4];
assign temp[1381] = ~window[28][5];
assign temp[1382] = window[28][6];
assign temp[1383] = window[28][7];
assign temp[1384] = ~window[28][8];
assign temp[1408] = window[29][0];
assign temp[1409] = window[29][1];
assign temp[1410] = window[29][2];
assign temp[1411] = ~window[29][3];
assign temp[1412] = ~window[29][4];
assign temp[1413] = ~window[29][5];
assign temp[1414] = ~window[29][6];
assign temp[1415] = window[29][7];
assign temp[1416] = window[29][8];
assign temp[1440] = window[30][0];
assign temp[1441] = ~window[30][1];
assign temp[1442] = window[30][2];
assign temp[1443] = window[30][3];
assign temp[1444] = ~window[30][4];
assign temp[1445] = ~window[30][5];
assign temp[1446] = window[30][6];
assign temp[1447] = ~window[30][7];
assign temp[1448] = window[30][8];
assign temp[1472] = ~window[31][0];
assign temp[1473] = window[31][1];
assign temp[1474] = window[31][2];
assign temp[1475] = ~window[31][3];
assign temp[1476] = ~window[31][4];
assign temp[1477] = ~window[31][5];
assign temp[1478] = window[31][6];
assign temp[1479] = window[31][7];
assign temp[1480] = ~window[31][8];
assign temp[512] = ~window[0][0];
assign temp[513] = ~window[0][1];
assign temp[514] = ~window[0][2];
assign temp[515] = ~window[0][3];
assign temp[516] = ~window[0][4];
assign temp[517] = ~window[0][5];
assign temp[518] = ~window[0][6];
assign temp[519] = ~window[0][7];
assign temp[520] = ~window[0][8];
assign temp[544] = ~window[1][0];
assign temp[545] = window[1][1];
assign temp[546] = window[1][2];
assign temp[547] = ~window[1][3];
assign temp[548] = ~window[1][4];
assign temp[549] = window[1][5];
assign temp[550] = window[1][6];
assign temp[551] = ~window[1][7];
assign temp[552] = window[1][8];
assign temp[576] = ~window[2][0];
assign temp[577] = ~window[2][1];
assign temp[578] = ~window[2][2];
assign temp[579] = ~window[2][3];
assign temp[580] = ~window[2][4];
assign temp[581] = ~window[2][5];
assign temp[582] = ~window[2][6];
assign temp[583] = window[2][7];
assign temp[584] = ~window[2][8];
assign temp[608] = window[3][0];
assign temp[609] = ~window[3][1];
assign temp[610] = window[3][2];
assign temp[611] = ~window[3][3];
assign temp[612] = ~window[3][4];
assign temp[613] = window[3][5];
assign temp[614] = ~window[3][6];
assign temp[615] = window[3][7];
assign temp[616] = ~window[3][8];
assign temp[640] = ~window[4][0];
assign temp[641] = ~window[4][1];
assign temp[642] = ~window[4][2];
assign temp[643] = window[4][3];
assign temp[644] = ~window[4][4];
assign temp[645] = ~window[4][5];
assign temp[646] = window[4][6];
assign temp[647] = ~window[4][7];
assign temp[648] = window[4][8];
assign temp[672] = ~window[5][0];
assign temp[673] = window[5][1];
assign temp[674] = window[5][2];
assign temp[675] = ~window[5][3];
assign temp[676] = window[5][4];
assign temp[677] = ~window[5][5];
assign temp[678] = window[5][6];
assign temp[679] = ~window[5][7];
assign temp[680] = ~window[5][8];
assign temp[704] = window[6][0];
assign temp[705] = ~window[6][1];
assign temp[706] = ~window[6][2];
assign temp[707] = ~window[6][3];
assign temp[708] = ~window[6][4];
assign temp[709] = ~window[6][5];
assign temp[710] = ~window[6][6];
assign temp[711] = ~window[6][7];
assign temp[712] = ~window[6][8];
assign temp[736] = ~window[7][0];
assign temp[737] = window[7][1];
assign temp[738] = window[7][2];
assign temp[739] = window[7][3];
assign temp[740] = window[7][4];
assign temp[741] = window[7][5];
assign temp[742] = window[7][6];
assign temp[743] = ~window[7][7];
assign temp[744] = window[7][8];
assign temp[768] = window[8][0];
assign temp[769] = ~window[8][1];
assign temp[770] = ~window[8][2];
assign temp[771] = ~window[8][3];
assign temp[772] = ~window[8][4];
assign temp[773] = ~window[8][5];
assign temp[774] = ~window[8][6];
assign temp[775] = ~window[8][7];
assign temp[776] = ~window[8][8];
assign temp[800] = window[9][0];
assign temp[801] = window[9][1];
assign temp[802] = window[9][2];
assign temp[803] = ~window[9][3];
assign temp[804] = window[9][4];
assign temp[805] = window[9][5];
assign temp[806] = ~window[9][6];
assign temp[807] = window[9][7];
assign temp[808] = window[9][8];
assign temp[832] = ~window[10][0];
assign temp[833] = window[10][1];
assign temp[834] = window[10][2];
assign temp[835] = window[10][3];
assign temp[836] = window[10][4];
assign temp[837] = window[10][5];
assign temp[838] = window[10][6];
assign temp[839] = window[10][7];
assign temp[840] = window[10][8];
assign temp[864] = ~window[11][0];
assign temp[865] = ~window[11][1];
assign temp[866] = ~window[11][2];
assign temp[867] = ~window[11][3];
assign temp[868] = ~window[11][4];
assign temp[869] = window[11][5];
assign temp[870] = window[11][6];
assign temp[871] = window[11][7];
assign temp[872] = window[11][8];
assign temp[896] = window[12][0];
assign temp[897] = ~window[12][1];
assign temp[898] = window[12][2];
assign temp[899] = ~window[12][3];
assign temp[900] = ~window[12][4];
assign temp[901] = ~window[12][5];
assign temp[902] = ~window[12][6];
assign temp[903] = window[12][7];
assign temp[904] = ~window[12][8];
assign temp[928] = ~window[13][0];
assign temp[929] = window[13][1];
assign temp[930] = window[13][2];
assign temp[931] = ~window[13][3];
assign temp[932] = window[13][4];
assign temp[933] = window[13][5];
assign temp[934] = ~window[13][6];
assign temp[935] = window[13][7];
assign temp[936] = ~window[13][8];
assign temp[960] = ~window[14][0];
assign temp[961] = window[14][1];
assign temp[962] = window[14][2];
assign temp[963] = window[14][3];
assign temp[964] = window[14][4];
assign temp[965] = ~window[14][5];
assign temp[966] = window[14][6];
assign temp[967] = window[14][7];
assign temp[968] = ~window[14][8];
assign temp[992] = window[15][0];
assign temp[993] = ~window[15][1];
assign temp[994] = ~window[15][2];
assign temp[995] = window[15][3];
assign temp[996] = ~window[15][4];
assign temp[997] = window[15][5];
assign temp[998] = window[15][6];
assign temp[999] = ~window[15][7];
assign temp[1000] = window[15][8];
assign temp[1024] = window[16][0];
assign temp[1025] = window[16][1];
assign temp[1026] = window[16][2];
assign temp[1027] = window[16][3];
assign temp[1028] = window[16][4];
assign temp[1029] = ~window[16][5];
assign temp[1030] = ~window[16][6];
assign temp[1031] = window[16][7];
assign temp[1032] = ~window[16][8];
assign temp[1056] = ~window[17][0];
assign temp[1057] = window[17][1];
assign temp[1058] = window[17][2];
assign temp[1059] = window[17][3];
assign temp[1060] = window[17][4];
assign temp[1061] = window[17][5];
assign temp[1062] = window[17][6];
assign temp[1063] = ~window[17][7];
assign temp[1064] = window[17][8];
assign temp[1088] = window[18][0];
assign temp[1089] = window[18][1];
assign temp[1090] = window[18][2];
assign temp[1091] = window[18][3];
assign temp[1092] = window[18][4];
assign temp[1093] = ~window[18][5];
assign temp[1094] = window[18][6];
assign temp[1095] = window[18][7];
assign temp[1096] = window[18][8];
assign temp[1120] = ~window[19][0];
assign temp[1121] = window[19][1];
assign temp[1122] = window[19][2];
assign temp[1123] = window[19][3];
assign temp[1124] = window[19][4];
assign temp[1125] = window[19][5];
assign temp[1126] = window[19][6];
assign temp[1127] = window[19][7];
assign temp[1128] = ~window[19][8];
assign temp[1152] = window[20][0];
assign temp[1153] = window[20][1];
assign temp[1154] = window[20][2];
assign temp[1155] = window[20][3];
assign temp[1156] = window[20][4];
assign temp[1157] = window[20][5];
assign temp[1158] = window[20][6];
assign temp[1159] = window[20][7];
assign temp[1160] = window[20][8];
assign temp[1184] = ~window[21][0];
assign temp[1185] = window[21][1];
assign temp[1186] = window[21][2];
assign temp[1187] = window[21][3];
assign temp[1188] = window[21][4];
assign temp[1189] = window[21][5];
assign temp[1190] = window[21][6];
assign temp[1191] = window[21][7];
assign temp[1192] = window[21][8];
assign temp[1216] = ~window[22][0];
assign temp[1217] = ~window[22][1];
assign temp[1218] = ~window[22][2];
assign temp[1219] = ~window[22][3];
assign temp[1220] = ~window[22][4];
assign temp[1221] = ~window[22][5];
assign temp[1222] = ~window[22][6];
assign temp[1223] = ~window[22][7];
assign temp[1224] = ~window[22][8];
assign temp[1248] = ~window[23][0];
assign temp[1249] = window[23][1];
assign temp[1250] = window[23][2];
assign temp[1251] = window[23][3];
assign temp[1252] = window[23][4];
assign temp[1253] = ~window[23][5];
assign temp[1254] = window[23][6];
assign temp[1255] = window[23][7];
assign temp[1256] = ~window[23][8];
assign temp[1280] = ~window[24][0];
assign temp[1281] = ~window[24][1];
assign temp[1282] = window[24][2];
assign temp[1283] = ~window[24][3];
assign temp[1284] = ~window[24][4];
assign temp[1285] = ~window[24][5];
assign temp[1286] = ~window[24][6];
assign temp[1287] = window[24][7];
assign temp[1288] = ~window[24][8];
assign temp[1312] = window[25][0];
assign temp[1313] = window[25][1];
assign temp[1314] = window[25][2];
assign temp[1315] = window[25][3];
assign temp[1316] = window[25][4];
assign temp[1317] = ~window[25][5];
assign temp[1318] = ~window[25][6];
assign temp[1319] = window[25][7];
assign temp[1320] = ~window[25][8];
assign temp[1344] = ~window[26][0];
assign temp[1345] = ~window[26][1];
assign temp[1346] = ~window[26][2];
assign temp[1347] = ~window[26][3];
assign temp[1348] = ~window[26][4];
assign temp[1349] = window[26][5];
assign temp[1350] = ~window[26][6];
assign temp[1351] = ~window[26][7];
assign temp[1352] = window[26][8];
assign temp[1376] = window[27][0];
assign temp[1377] = window[27][1];
assign temp[1378] = window[27][2];
assign temp[1379] = window[27][3];
assign temp[1380] = window[27][4];
assign temp[1381] = window[27][5];
assign temp[1382] = window[27][6];
assign temp[1383] = window[27][7];
assign temp[1384] = window[27][8];
assign temp[1408] = ~window[28][0];
assign temp[1409] = ~window[28][1];
assign temp[1410] = window[28][2];
assign temp[1411] = ~window[28][3];
assign temp[1412] = window[28][4];
assign temp[1413] = window[28][5];
assign temp[1414] = window[28][6];
assign temp[1415] = window[28][7];
assign temp[1416] = window[28][8];
assign temp[1440] = ~window[29][0];
assign temp[1441] = ~window[29][1];
assign temp[1442] = ~window[29][2];
assign temp[1443] = ~window[29][3];
assign temp[1444] = window[29][4];
assign temp[1445] = ~window[29][5];
assign temp[1446] = window[29][6];
assign temp[1447] = ~window[29][7];
assign temp[1448] = ~window[29][8];
assign temp[1472] = ~window[30][0];
assign temp[1473] = window[30][1];
assign temp[1474] = window[30][2];
assign temp[1475] = window[30][3];
assign temp[1476] = window[30][4];
assign temp[1477] = ~window[30][5];
assign temp[1478] = ~window[30][6];
assign temp[1479] = ~window[30][7];
assign temp[1480] = ~window[30][8];
assign temp[1504] = ~window[31][0];
assign temp[1505] = ~window[31][1];
assign temp[1506] = window[31][2];
assign temp[1507] = ~window[31][3];
assign temp[1508] = ~window[31][4];
assign temp[1509] = ~window[31][5];
assign temp[1510] = ~window[31][6];
assign temp[1511] = ~window[31][7];
assign temp[1512] = ~window[31][8];
assign temp[544] = ~window[0][0];
assign temp[545] = ~window[0][1];
assign temp[546] = window[0][2];
assign temp[547] = window[0][3];
assign temp[548] = window[0][4];
assign temp[549] = ~window[0][5];
assign temp[550] = window[0][6];
assign temp[551] = window[0][7];
assign temp[552] = window[0][8];
assign temp[576] = window[1][0];
assign temp[577] = window[1][1];
assign temp[578] = window[1][2];
assign temp[579] = window[1][3];
assign temp[580] = window[1][4];
assign temp[581] = ~window[1][5];
assign temp[582] = window[1][6];
assign temp[583] = window[1][7];
assign temp[584] = ~window[1][8];
assign temp[608] = ~window[2][0];
assign temp[609] = ~window[2][1];
assign temp[610] = window[2][2];
assign temp[611] = window[2][3];
assign temp[612] = window[2][4];
assign temp[613] = window[2][5];
assign temp[614] = window[2][6];
assign temp[615] = ~window[2][7];
assign temp[616] = ~window[2][8];
assign temp[640] = window[3][0];
assign temp[641] = ~window[3][1];
assign temp[642] = window[3][2];
assign temp[643] = window[3][3];
assign temp[644] = window[3][4];
assign temp[645] = window[3][5];
assign temp[646] = ~window[3][6];
assign temp[647] = ~window[3][7];
assign temp[648] = ~window[3][8];
assign temp[672] = ~window[4][0];
assign temp[673] = ~window[4][1];
assign temp[674] = ~window[4][2];
assign temp[675] = window[4][3];
assign temp[676] = ~window[4][4];
assign temp[677] = ~window[4][5];
assign temp[678] = window[4][6];
assign temp[679] = window[4][7];
assign temp[680] = window[4][8];
assign temp[704] = window[5][0];
assign temp[705] = window[5][1];
assign temp[706] = window[5][2];
assign temp[707] = ~window[5][3];
assign temp[708] = ~window[5][4];
assign temp[709] = window[5][5];
assign temp[710] = window[5][6];
assign temp[711] = window[5][7];
assign temp[712] = window[5][8];
assign temp[736] = ~window[6][0];
assign temp[737] = ~window[6][1];
assign temp[738] = ~window[6][2];
assign temp[739] = ~window[6][3];
assign temp[740] = window[6][4];
assign temp[741] = ~window[6][5];
assign temp[742] = ~window[6][6];
assign temp[743] = window[6][7];
assign temp[744] = ~window[6][8];
assign temp[768] = window[7][0];
assign temp[769] = ~window[7][1];
assign temp[770] = ~window[7][2];
assign temp[771] = window[7][3];
assign temp[772] = ~window[7][4];
assign temp[773] = ~window[7][5];
assign temp[774] = window[7][6];
assign temp[775] = window[7][7];
assign temp[776] = window[7][8];
assign temp[800] = ~window[8][0];
assign temp[801] = window[8][1];
assign temp[802] = window[8][2];
assign temp[803] = window[8][3];
assign temp[804] = ~window[8][4];
assign temp[805] = ~window[8][5];
assign temp[806] = window[8][6];
assign temp[807] = window[8][7];
assign temp[808] = window[8][8];
assign temp[832] = window[9][0];
assign temp[833] = window[9][1];
assign temp[834] = window[9][2];
assign temp[835] = window[9][3];
assign temp[836] = window[9][4];
assign temp[837] = window[9][5];
assign temp[838] = window[9][6];
assign temp[839] = ~window[9][7];
assign temp[840] = ~window[9][8];
assign temp[864] = ~window[10][0];
assign temp[865] = window[10][1];
assign temp[866] = ~window[10][2];
assign temp[867] = window[10][3];
assign temp[868] = window[10][4];
assign temp[869] = ~window[10][5];
assign temp[870] = window[10][6];
assign temp[871] = window[10][7];
assign temp[872] = ~window[10][8];
assign temp[896] = ~window[11][0];
assign temp[897] = ~window[11][1];
assign temp[898] = ~window[11][2];
assign temp[899] = ~window[11][3];
assign temp[900] = window[11][4];
assign temp[901] = window[11][5];
assign temp[902] = window[11][6];
assign temp[903] = window[11][7];
assign temp[904] = window[11][8];
assign temp[928] = window[12][0];
assign temp[929] = window[12][1];
assign temp[930] = window[12][2];
assign temp[931] = window[12][3];
assign temp[932] = window[12][4];
assign temp[933] = window[12][5];
assign temp[934] = ~window[12][6];
assign temp[935] = window[12][7];
assign temp[936] = window[12][8];
assign temp[960] = window[13][0];
assign temp[961] = window[13][1];
assign temp[962] = window[13][2];
assign temp[963] = window[13][3];
assign temp[964] = window[13][4];
assign temp[965] = window[13][5];
assign temp[966] = window[13][6];
assign temp[967] = window[13][7];
assign temp[968] = window[13][8];
assign temp[992] = ~window[14][0];
assign temp[993] = ~window[14][1];
assign temp[994] = window[14][2];
assign temp[995] = window[14][3];
assign temp[996] = ~window[14][4];
assign temp[997] = ~window[14][5];
assign temp[998] = window[14][6];
assign temp[999] = window[14][7];
assign temp[1000] = window[14][8];
assign temp[1024] = window[15][0];
assign temp[1025] = ~window[15][1];
assign temp[1026] = ~window[15][2];
assign temp[1027] = ~window[15][3];
assign temp[1028] = window[15][4];
assign temp[1029] = window[15][5];
assign temp[1030] = window[15][6];
assign temp[1031] = ~window[15][7];
assign temp[1032] = ~window[15][8];
assign temp[1056] = window[16][0];
assign temp[1057] = window[16][1];
assign temp[1058] = ~window[16][2];
assign temp[1059] = ~window[16][3];
assign temp[1060] = ~window[16][4];
assign temp[1061] = window[16][5];
assign temp[1062] = window[16][6];
assign temp[1063] = window[16][7];
assign temp[1064] = window[16][8];
assign temp[1088] = window[17][0];
assign temp[1089] = window[17][1];
assign temp[1090] = window[17][2];
assign temp[1091] = window[17][3];
assign temp[1092] = window[17][4];
assign temp[1093] = ~window[17][5];
assign temp[1094] = window[17][6];
assign temp[1095] = ~window[17][7];
assign temp[1096] = ~window[17][8];
assign temp[1120] = window[18][0];
assign temp[1121] = window[18][1];
assign temp[1122] = ~window[18][2];
assign temp[1123] = window[18][3];
assign temp[1124] = window[18][4];
assign temp[1125] = ~window[18][5];
assign temp[1126] = ~window[18][6];
assign temp[1127] = ~window[18][7];
assign temp[1128] = window[18][8];
assign temp[1152] = ~window[19][0];
assign temp[1153] = ~window[19][1];
assign temp[1154] = ~window[19][2];
assign temp[1155] = window[19][3];
assign temp[1156] = window[19][4];
assign temp[1157] = window[19][5];
assign temp[1158] = ~window[19][6];
assign temp[1159] = window[19][7];
assign temp[1160] = ~window[19][8];
assign temp[1184] = window[20][0];
assign temp[1185] = window[20][1];
assign temp[1186] = window[20][2];
assign temp[1187] = window[20][3];
assign temp[1188] = window[20][4];
assign temp[1189] = window[20][5];
assign temp[1190] = ~window[20][6];
assign temp[1191] = ~window[20][7];
assign temp[1192] = ~window[20][8];
assign temp[1216] = ~window[21][0];
assign temp[1217] = ~window[21][1];
assign temp[1218] = ~window[21][2];
assign temp[1219] = ~window[21][3];
assign temp[1220] = window[21][4];
assign temp[1221] = ~window[21][5];
assign temp[1222] = window[21][6];
assign temp[1223] = window[21][7];
assign temp[1224] = ~window[21][8];
assign temp[1248] = window[22][0];
assign temp[1249] = ~window[22][1];
assign temp[1250] = ~window[22][2];
assign temp[1251] = window[22][3];
assign temp[1252] = ~window[22][4];
assign temp[1253] = ~window[22][5];
assign temp[1254] = window[22][6];
assign temp[1255] = window[22][7];
assign temp[1256] = window[22][8];
assign temp[1280] = ~window[23][0];
assign temp[1281] = window[23][1];
assign temp[1282] = window[23][2];
assign temp[1283] = window[23][3];
assign temp[1284] = ~window[23][4];
assign temp[1285] = ~window[23][5];
assign temp[1286] = window[23][6];
assign temp[1287] = ~window[23][7];
assign temp[1288] = window[23][8];
assign temp[1312] = ~window[24][0];
assign temp[1313] = window[24][1];
assign temp[1314] = window[24][2];
assign temp[1315] = ~window[24][3];
assign temp[1316] = window[24][4];
assign temp[1317] = window[24][5];
assign temp[1318] = window[24][6];
assign temp[1319] = ~window[24][7];
assign temp[1320] = window[24][8];
assign temp[1344] = ~window[25][0];
assign temp[1345] = window[25][1];
assign temp[1346] = window[25][2];
assign temp[1347] = ~window[25][3];
assign temp[1348] = ~window[25][4];
assign temp[1349] = ~window[25][5];
assign temp[1350] = window[25][6];
assign temp[1351] = window[25][7];
assign temp[1352] = window[25][8];
assign temp[1376] = window[26][0];
assign temp[1377] = ~window[26][1];
assign temp[1378] = ~window[26][2];
assign temp[1379] = window[26][3];
assign temp[1380] = window[26][4];
assign temp[1381] = ~window[26][5];
assign temp[1382] = window[26][6];
assign temp[1383] = window[26][7];
assign temp[1384] = ~window[26][8];
assign temp[1408] = window[27][0];
assign temp[1409] = ~window[27][1];
assign temp[1410] = ~window[27][2];
assign temp[1411] = window[27][3];
assign temp[1412] = ~window[27][4];
assign temp[1413] = ~window[27][5];
assign temp[1414] = window[27][6];
assign temp[1415] = ~window[27][7];
assign temp[1416] = window[27][8];
assign temp[1440] = window[28][0];
assign temp[1441] = window[28][1];
assign temp[1442] = ~window[28][2];
assign temp[1443] = ~window[28][3];
assign temp[1444] = window[28][4];
assign temp[1445] = window[28][5];
assign temp[1446] = window[28][6];
assign temp[1447] = window[28][7];
assign temp[1448] = window[28][8];
assign temp[1472] = window[29][0];
assign temp[1473] = window[29][1];
assign temp[1474] = ~window[29][2];
assign temp[1475] = window[29][3];
assign temp[1476] = window[29][4];
assign temp[1477] = ~window[29][5];
assign temp[1478] = window[29][6];
assign temp[1479] = window[29][7];
assign temp[1480] = window[29][8];
assign temp[1504] = window[30][0];
assign temp[1505] = window[30][1];
assign temp[1506] = window[30][2];
assign temp[1507] = window[30][3];
assign temp[1508] = ~window[30][4];
assign temp[1509] = ~window[30][5];
assign temp[1510] = ~window[30][6];
assign temp[1511] = window[30][7];
assign temp[1512] = window[30][8];
assign temp[1536] = ~window[31][0];
assign temp[1537] = window[31][1];
assign temp[1538] = window[31][2];
assign temp[1539] = window[31][3];
assign temp[1540] = window[31][4];
assign temp[1541] = window[31][5];
assign temp[1542] = window[31][6];
assign temp[1543] = ~window[31][7];
assign temp[1544] = window[31][8];
assign temp[576] = ~window[0][0];
assign temp[577] = ~window[0][1];
assign temp[578] = ~window[0][2];
assign temp[579] = window[0][3];
assign temp[580] = window[0][4];
assign temp[581] = window[0][5];
assign temp[582] = ~window[0][6];
assign temp[583] = window[0][7];
assign temp[584] = ~window[0][8];
assign temp[608] = window[1][0];
assign temp[609] = window[1][1];
assign temp[610] = ~window[1][2];
assign temp[611] = ~window[1][3];
assign temp[612] = window[1][4];
assign temp[613] = window[1][5];
assign temp[614] = window[1][6];
assign temp[615] = window[1][7];
assign temp[616] = window[1][8];
assign temp[640] = ~window[2][0];
assign temp[641] = ~window[2][1];
assign temp[642] = ~window[2][2];
assign temp[643] = window[2][3];
assign temp[644] = window[2][4];
assign temp[645] = window[2][5];
assign temp[646] = window[2][6];
assign temp[647] = window[2][7];
assign temp[648] = ~window[2][8];
assign temp[672] = ~window[3][0];
assign temp[673] = ~window[3][1];
assign temp[674] = ~window[3][2];
assign temp[675] = window[3][3];
assign temp[676] = window[3][4];
assign temp[677] = window[3][5];
assign temp[678] = window[3][6];
assign temp[679] = ~window[3][7];
assign temp[680] = ~window[3][8];
assign temp[704] = ~window[4][0];
assign temp[705] = ~window[4][1];
assign temp[706] = window[4][2];
assign temp[707] = ~window[4][3];
assign temp[708] = ~window[4][4];
assign temp[709] = ~window[4][5];
assign temp[710] = ~window[4][6];
assign temp[711] = ~window[4][7];
assign temp[712] = ~window[4][8];
assign temp[736] = window[5][0];
assign temp[737] = ~window[5][1];
assign temp[738] = ~window[5][2];
assign temp[739] = window[5][3];
assign temp[740] = window[5][4];
assign temp[741] = ~window[5][5];
assign temp[742] = ~window[5][6];
assign temp[743] = ~window[5][7];
assign temp[744] = ~window[5][8];
assign temp[768] = ~window[6][0];
assign temp[769] = ~window[6][1];
assign temp[770] = ~window[6][2];
assign temp[771] = window[6][3];
assign temp[772] = ~window[6][4];
assign temp[773] = window[6][5];
assign temp[774] = window[6][6];
assign temp[775] = window[6][7];
assign temp[776] = ~window[6][8];
assign temp[800] = window[7][0];
assign temp[801] = ~window[7][1];
assign temp[802] = window[7][2];
assign temp[803] = window[7][3];
assign temp[804] = window[7][4];
assign temp[805] = ~window[7][5];
assign temp[806] = ~window[7][6];
assign temp[807] = ~window[7][7];
assign temp[808] = ~window[7][8];
assign temp[832] = ~window[8][0];
assign temp[833] = window[8][1];
assign temp[834] = window[8][2];
assign temp[835] = window[8][3];
assign temp[836] = window[8][4];
assign temp[837] = window[8][5];
assign temp[838] = window[8][6];
assign temp[839] = ~window[8][7];
assign temp[840] = ~window[8][8];
assign temp[864] = window[9][0];
assign temp[865] = ~window[9][1];
assign temp[866] = ~window[9][2];
assign temp[867] = window[9][3];
assign temp[868] = window[9][4];
assign temp[869] = window[9][5];
assign temp[870] = window[9][6];
assign temp[871] = window[9][7];
assign temp[872] = ~window[9][8];
assign temp[896] = window[10][0];
assign temp[897] = ~window[10][1];
assign temp[898] = ~window[10][2];
assign temp[899] = window[10][3];
assign temp[900] = window[10][4];
assign temp[901] = window[10][5];
assign temp[902] = ~window[10][6];
assign temp[903] = ~window[10][7];
assign temp[904] = ~window[10][8];
assign temp[928] = window[11][0];
assign temp[929] = window[11][1];
assign temp[930] = window[11][2];
assign temp[931] = window[11][3];
assign temp[932] = window[11][4];
assign temp[933] = ~window[11][5];
assign temp[934] = ~window[11][6];
assign temp[935] = ~window[11][7];
assign temp[936] = window[11][8];
assign temp[960] = ~window[12][0];
assign temp[961] = window[12][1];
assign temp[962] = ~window[12][2];
assign temp[963] = ~window[12][3];
assign temp[964] = ~window[12][4];
assign temp[965] = window[12][5];
assign temp[966] = window[12][6];
assign temp[967] = window[12][7];
assign temp[968] = window[12][8];
assign temp[992] = ~window[13][0];
assign temp[993] = window[13][1];
assign temp[994] = window[13][2];
assign temp[995] = ~window[13][3];
assign temp[996] = ~window[13][4];
assign temp[997] = ~window[13][5];
assign temp[998] = ~window[13][6];
assign temp[999] = window[13][7];
assign temp[1000] = window[13][8];
assign temp[1024] = ~window[14][0];
assign temp[1025] = ~window[14][1];
assign temp[1026] = window[14][2];
assign temp[1027] = window[14][3];
assign temp[1028] = window[14][4];
assign temp[1029] = ~window[14][5];
assign temp[1030] = ~window[14][6];
assign temp[1031] = ~window[14][7];
assign temp[1032] = ~window[14][8];
assign temp[1056] = ~window[15][0];
assign temp[1057] = window[15][1];
assign temp[1058] = window[15][2];
assign temp[1059] = window[15][3];
assign temp[1060] = ~window[15][4];
assign temp[1061] = ~window[15][5];
assign temp[1062] = ~window[15][6];
assign temp[1063] = window[15][7];
assign temp[1064] = ~window[15][8];
assign temp[1088] = ~window[16][0];
assign temp[1089] = window[16][1];
assign temp[1090] = window[16][2];
assign temp[1091] = window[16][3];
assign temp[1092] = window[16][4];
assign temp[1093] = ~window[16][5];
assign temp[1094] = ~window[16][6];
assign temp[1095] = ~window[16][7];
assign temp[1096] = ~window[16][8];
assign temp[1120] = window[17][0];
assign temp[1121] = ~window[17][1];
assign temp[1122] = ~window[17][2];
assign temp[1123] = ~window[17][3];
assign temp[1124] = window[17][4];
assign temp[1125] = window[17][5];
assign temp[1126] = window[17][6];
assign temp[1127] = window[17][7];
assign temp[1128] = ~window[17][8];
assign temp[1152] = window[18][0];
assign temp[1153] = window[18][1];
assign temp[1154] = ~window[18][2];
assign temp[1155] = ~window[18][3];
assign temp[1156] = ~window[18][4];
assign temp[1157] = window[18][5];
assign temp[1158] = ~window[18][6];
assign temp[1159] = ~window[18][7];
assign temp[1160] = ~window[18][8];
assign temp[1184] = window[19][0];
assign temp[1185] = ~window[19][1];
assign temp[1186] = ~window[19][2];
assign temp[1187] = ~window[19][3];
assign temp[1188] = ~window[19][4];
assign temp[1189] = ~window[19][5];
assign temp[1190] = ~window[19][6];
assign temp[1191] = window[19][7];
assign temp[1192] = window[19][8];
assign temp[1216] = ~window[20][0];
assign temp[1217] = window[20][1];
assign temp[1218] = ~window[20][2];
assign temp[1219] = ~window[20][3];
assign temp[1220] = window[20][4];
assign temp[1221] = window[20][5];
assign temp[1222] = window[20][6];
assign temp[1223] = window[20][7];
assign temp[1224] = ~window[20][8];
assign temp[1248] = window[21][0];
assign temp[1249] = ~window[21][1];
assign temp[1250] = ~window[21][2];
assign temp[1251] = window[21][3];
assign temp[1252] = ~window[21][4];
assign temp[1253] = ~window[21][5];
assign temp[1254] = ~window[21][6];
assign temp[1255] = ~window[21][7];
assign temp[1256] = ~window[21][8];
assign temp[1280] = window[22][0];
assign temp[1281] = window[22][1];
assign temp[1282] = window[22][2];
assign temp[1283] = ~window[22][3];
assign temp[1284] = window[22][4];
assign temp[1285] = ~window[22][5];
assign temp[1286] = ~window[22][6];
assign temp[1287] = window[22][7];
assign temp[1288] = window[22][8];
assign temp[1312] = ~window[23][0];
assign temp[1313] = ~window[23][1];
assign temp[1314] = ~window[23][2];
assign temp[1315] = window[23][3];
assign temp[1316] = window[23][4];
assign temp[1317] = window[23][5];
assign temp[1318] = window[23][6];
assign temp[1319] = ~window[23][7];
assign temp[1320] = ~window[23][8];
assign temp[1344] = ~window[24][0];
assign temp[1345] = ~window[24][1];
assign temp[1346] = ~window[24][2];
assign temp[1347] = window[24][3];
assign temp[1348] = ~window[24][4];
assign temp[1349] = ~window[24][5];
assign temp[1350] = window[24][6];
assign temp[1351] = window[24][7];
assign temp[1352] = ~window[24][8];
assign temp[1376] = ~window[25][0];
assign temp[1377] = ~window[25][1];
assign temp[1378] = window[25][2];
assign temp[1379] = ~window[25][3];
assign temp[1380] = window[25][4];
assign temp[1381] = ~window[25][5];
assign temp[1382] = window[25][6];
assign temp[1383] = ~window[25][7];
assign temp[1384] = ~window[25][8];
assign temp[1408] = ~window[26][0];
assign temp[1409] = ~window[26][1];
assign temp[1410] = ~window[26][2];
assign temp[1411] = window[26][3];
assign temp[1412] = ~window[26][4];
assign temp[1413] = window[26][5];
assign temp[1414] = ~window[26][6];
assign temp[1415] = window[26][7];
assign temp[1416] = window[26][8];
assign temp[1440] = ~window[27][0];
assign temp[1441] = window[27][1];
assign temp[1442] = window[27][2];
assign temp[1443] = ~window[27][3];
assign temp[1444] = window[27][4];
assign temp[1445] = ~window[27][5];
assign temp[1446] = ~window[27][6];
assign temp[1447] = ~window[27][7];
assign temp[1448] = ~window[27][8];
assign temp[1472] = ~window[28][0];
assign temp[1473] = window[28][1];
assign temp[1474] = window[28][2];
assign temp[1475] = ~window[28][3];
assign temp[1476] = ~window[28][4];
assign temp[1477] = ~window[28][5];
assign temp[1478] = ~window[28][6];
assign temp[1479] = window[28][7];
assign temp[1480] = ~window[28][8];
assign temp[1504] = window[29][0];
assign temp[1505] = window[29][1];
assign temp[1506] = window[29][2];
assign temp[1507] = ~window[29][3];
assign temp[1508] = window[29][4];
assign temp[1509] = ~window[29][5];
assign temp[1510] = ~window[29][6];
assign temp[1511] = ~window[29][7];
assign temp[1512] = window[29][8];
assign temp[1536] = window[30][0];
assign temp[1537] = window[30][1];
assign temp[1538] = window[30][2];
assign temp[1539] = ~window[30][3];
assign temp[1540] = ~window[30][4];
assign temp[1541] = ~window[30][5];
assign temp[1542] = ~window[30][6];
assign temp[1543] = ~window[30][7];
assign temp[1544] = window[30][8];
assign temp[1568] = ~window[31][0];
assign temp[1569] = ~window[31][1];
assign temp[1570] = ~window[31][2];
assign temp[1571] = window[31][3];
assign temp[1572] = window[31][4];
assign temp[1573] = ~window[31][5];
assign temp[1574] = window[31][6];
assign temp[1575] = window[31][7];
assign temp[1576] = window[31][8];
assign temp[608] = window[0][0];
assign temp[609] = ~window[0][1];
assign temp[610] = window[0][2];
assign temp[611] = window[0][3];
assign temp[612] = ~window[0][4];
assign temp[613] = window[0][5];
assign temp[614] = window[0][6];
assign temp[615] = ~window[0][7];
assign temp[616] = ~window[0][8];
assign temp[640] = window[1][0];
assign temp[641] = ~window[1][1];
assign temp[642] = ~window[1][2];
assign temp[643] = window[1][3];
assign temp[644] = window[1][4];
assign temp[645] = ~window[1][5];
assign temp[646] = window[1][6];
assign temp[647] = window[1][7];
assign temp[648] = window[1][8];
assign temp[672] = window[2][0];
assign temp[673] = ~window[2][1];
assign temp[674] = ~window[2][2];
assign temp[675] = ~window[2][3];
assign temp[676] = window[2][4];
assign temp[677] = window[2][5];
assign temp[678] = ~window[2][6];
assign temp[679] = ~window[2][7];
assign temp[680] = window[2][8];
assign temp[704] = window[3][0];
assign temp[705] = window[3][1];
assign temp[706] = window[3][2];
assign temp[707] = ~window[3][3];
assign temp[708] = window[3][4];
assign temp[709] = window[3][5];
assign temp[710] = ~window[3][6];
assign temp[711] = ~window[3][7];
assign temp[712] = window[3][8];
assign temp[736] = ~window[4][0];
assign temp[737] = window[4][1];
assign temp[738] = window[4][2];
assign temp[739] = window[4][3];
assign temp[740] = window[4][4];
assign temp[741] = window[4][5];
assign temp[742] = window[4][6];
assign temp[743] = window[4][7];
assign temp[744] = ~window[4][8];
assign temp[768] = window[5][0];
assign temp[769] = ~window[5][1];
assign temp[770] = ~window[5][2];
assign temp[771] = ~window[5][3];
assign temp[772] = ~window[5][4];
assign temp[773] = ~window[5][5];
assign temp[774] = window[5][6];
assign temp[775] = ~window[5][7];
assign temp[776] = ~window[5][8];
assign temp[800] = window[6][0];
assign temp[801] = ~window[6][1];
assign temp[802] = ~window[6][2];
assign temp[803] = ~window[6][3];
assign temp[804] = window[6][4];
assign temp[805] = ~window[6][5];
assign temp[806] = ~window[6][6];
assign temp[807] = ~window[6][7];
assign temp[808] = window[6][8];
assign temp[832] = ~window[7][0];
assign temp[833] = window[7][1];
assign temp[834] = ~window[7][2];
assign temp[835] = window[7][3];
assign temp[836] = window[7][4];
assign temp[837] = window[7][5];
assign temp[838] = window[7][6];
assign temp[839] = window[7][7];
assign temp[840] = ~window[7][8];
assign temp[864] = window[8][0];
assign temp[865] = window[8][1];
assign temp[866] = window[8][2];
assign temp[867] = window[8][3];
assign temp[868] = window[8][4];
assign temp[869] = window[8][5];
assign temp[870] = window[8][6];
assign temp[871] = window[8][7];
assign temp[872] = window[8][8];
assign temp[896] = window[9][0];
assign temp[897] = window[9][1];
assign temp[898] = ~window[9][2];
assign temp[899] = window[9][3];
assign temp[900] = window[9][4];
assign temp[901] = window[9][5];
assign temp[902] = ~window[9][6];
assign temp[903] = window[9][7];
assign temp[904] = window[9][8];
assign temp[928] = window[10][0];
assign temp[929] = window[10][1];
assign temp[930] = ~window[10][2];
assign temp[931] = window[10][3];
assign temp[932] = window[10][4];
assign temp[933] = window[10][5];
assign temp[934] = window[10][6];
assign temp[935] = window[10][7];
assign temp[936] = window[10][8];
assign temp[960] = ~window[11][0];
assign temp[961] = window[11][1];
assign temp[962] = window[11][2];
assign temp[963] = ~window[11][3];
assign temp[964] = window[11][4];
assign temp[965] = ~window[11][5];
assign temp[966] = window[11][6];
assign temp[967] = ~window[11][7];
assign temp[968] = ~window[11][8];
assign temp[992] = ~window[12][0];
assign temp[993] = ~window[12][1];
assign temp[994] = window[12][2];
assign temp[995] = window[12][3];
assign temp[996] = window[12][4];
assign temp[997] = window[12][5];
assign temp[998] = window[12][6];
assign temp[999] = window[12][7];
assign temp[1000] = window[12][8];
assign temp[1024] = window[13][0];
assign temp[1025] = window[13][1];
assign temp[1026] = window[13][2];
assign temp[1027] = window[13][3];
assign temp[1028] = window[13][4];
assign temp[1029] = window[13][5];
assign temp[1030] = window[13][6];
assign temp[1031] = window[13][7];
assign temp[1032] = ~window[13][8];
assign temp[1056] = ~window[14][0];
assign temp[1057] = ~window[14][1];
assign temp[1058] = ~window[14][2];
assign temp[1059] = window[14][3];
assign temp[1060] = window[14][4];
assign temp[1061] = window[14][5];
assign temp[1062] = window[14][6];
assign temp[1063] = window[14][7];
assign temp[1064] = window[14][8];
assign temp[1088] = ~window[15][0];
assign temp[1089] = window[15][1];
assign temp[1090] = ~window[15][2];
assign temp[1091] = window[15][3];
assign temp[1092] = window[15][4];
assign temp[1093] = window[15][5];
assign temp[1094] = window[15][6];
assign temp[1095] = window[15][7];
assign temp[1096] = window[15][8];
assign temp[1120] = window[16][0];
assign temp[1121] = window[16][1];
assign temp[1122] = window[16][2];
assign temp[1123] = window[16][3];
assign temp[1124] = window[16][4];
assign temp[1125] = window[16][5];
assign temp[1126] = window[16][6];
assign temp[1127] = window[16][7];
assign temp[1128] = ~window[16][8];
assign temp[1152] = ~window[17][0];
assign temp[1153] = ~window[17][1];
assign temp[1154] = window[17][2];
assign temp[1155] = ~window[17][3];
assign temp[1156] = window[17][4];
assign temp[1157] = ~window[17][5];
assign temp[1158] = window[17][6];
assign temp[1159] = window[17][7];
assign temp[1160] = window[17][8];
assign temp[1184] = window[18][0];
assign temp[1185] = window[18][1];
assign temp[1186] = window[18][2];
assign temp[1187] = window[18][3];
assign temp[1188] = window[18][4];
assign temp[1189] = window[18][5];
assign temp[1190] = ~window[18][6];
assign temp[1191] = window[18][7];
assign temp[1192] = window[18][8];
assign temp[1216] = window[19][0];
assign temp[1217] = ~window[19][1];
assign temp[1218] = window[19][2];
assign temp[1219] = ~window[19][3];
assign temp[1220] = ~window[19][4];
assign temp[1221] = ~window[19][5];
assign temp[1222] = window[19][6];
assign temp[1223] = ~window[19][7];
assign temp[1224] = ~window[19][8];
assign temp[1248] = window[20][0];
assign temp[1249] = window[20][1];
assign temp[1250] = window[20][2];
assign temp[1251] = ~window[20][3];
assign temp[1252] = window[20][4];
assign temp[1253] = window[20][5];
assign temp[1254] = ~window[20][6];
assign temp[1255] = window[20][7];
assign temp[1256] = window[20][8];
assign temp[1280] = window[21][0];
assign temp[1281] = window[21][1];
assign temp[1282] = ~window[21][2];
assign temp[1283] = window[21][3];
assign temp[1284] = ~window[21][4];
assign temp[1285] = ~window[21][5];
assign temp[1286] = window[21][6];
assign temp[1287] = window[21][7];
assign temp[1288] = ~window[21][8];
assign temp[1312] = ~window[22][0];
assign temp[1313] = ~window[22][1];
assign temp[1314] = window[22][2];
assign temp[1315] = window[22][3];
assign temp[1316] = ~window[22][4];
assign temp[1317] = window[22][5];
assign temp[1318] = window[22][6];
assign temp[1319] = window[22][7];
assign temp[1320] = window[22][8];
assign temp[1344] = window[23][0];
assign temp[1345] = ~window[23][1];
assign temp[1346] = ~window[23][2];
assign temp[1347] = window[23][3];
assign temp[1348] = ~window[23][4];
assign temp[1349] = window[23][5];
assign temp[1350] = window[23][6];
assign temp[1351] = ~window[23][7];
assign temp[1352] = window[23][8];
assign temp[1376] = window[24][0];
assign temp[1377] = window[24][1];
assign temp[1378] = window[24][2];
assign temp[1379] = window[24][3];
assign temp[1380] = window[24][4];
assign temp[1381] = window[24][5];
assign temp[1382] = ~window[24][6];
assign temp[1383] = ~window[24][7];
assign temp[1384] = window[24][8];
assign temp[1408] = ~window[25][0];
assign temp[1409] = window[25][1];
assign temp[1410] = ~window[25][2];
assign temp[1411] = window[25][3];
assign temp[1412] = window[25][4];
assign temp[1413] = window[25][5];
assign temp[1414] = window[25][6];
assign temp[1415] = ~window[25][7];
assign temp[1416] = window[25][8];
assign temp[1440] = window[26][0];
assign temp[1441] = ~window[26][1];
assign temp[1442] = ~window[26][2];
assign temp[1443] = ~window[26][3];
assign temp[1444] = ~window[26][4];
assign temp[1445] = ~window[26][5];
assign temp[1446] = window[26][6];
assign temp[1447] = window[26][7];
assign temp[1448] = ~window[26][8];
assign temp[1472] = ~window[27][0];
assign temp[1473] = window[27][1];
assign temp[1474] = window[27][2];
assign temp[1475] = window[27][3];
assign temp[1476] = window[27][4];
assign temp[1477] = window[27][5];
assign temp[1478] = window[27][6];
assign temp[1479] = window[27][7];
assign temp[1480] = ~window[27][8];
assign temp[1504] = window[28][0];
assign temp[1505] = window[28][1];
assign temp[1506] = window[28][2];
assign temp[1507] = window[28][3];
assign temp[1508] = window[28][4];
assign temp[1509] = window[28][5];
assign temp[1510] = window[28][6];
assign temp[1511] = window[28][7];
assign temp[1512] = window[28][8];
assign temp[1536] = ~window[29][0];
assign temp[1537] = ~window[29][1];
assign temp[1538] = window[29][2];
assign temp[1539] = ~window[29][3];
assign temp[1540] = ~window[29][4];
assign temp[1541] = window[29][5];
assign temp[1542] = window[29][6];
assign temp[1543] = window[29][7];
assign temp[1544] = ~window[29][8];
assign temp[1568] = ~window[30][0];
assign temp[1569] = ~window[30][1];
assign temp[1570] = window[30][2];
assign temp[1571] = window[30][3];
assign temp[1572] = ~window[30][4];
assign temp[1573] = ~window[30][5];
assign temp[1574] = window[30][6];
assign temp[1575] = ~window[30][7];
assign temp[1576] = ~window[30][8];
assign temp[1600] = ~window[31][0];
assign temp[1601] = ~window[31][1];
assign temp[1602] = ~window[31][2];
assign temp[1603] = window[31][3];
assign temp[1604] = window[31][4];
assign temp[1605] = window[31][5];
assign temp[1606] = window[31][6];
assign temp[1607] = window[31][7];
assign temp[1608] = window[31][8];
assign temp[640] = window[0][0];
assign temp[641] = window[0][1];
assign temp[642] = ~window[0][2];
assign temp[643] = window[0][3];
assign temp[644] = ~window[0][4];
assign temp[645] = ~window[0][5];
assign temp[646] = window[0][6];
assign temp[647] = ~window[0][7];
assign temp[648] = ~window[0][8];
assign temp[672] = window[1][0];
assign temp[673] = window[1][1];
assign temp[674] = ~window[1][2];
assign temp[675] = window[1][3];
assign temp[676] = window[1][4];
assign temp[677] = window[1][5];
assign temp[678] = window[1][6];
assign temp[679] = ~window[1][7];
assign temp[680] = ~window[1][8];
assign temp[704] = window[2][0];
assign temp[705] = ~window[2][1];
assign temp[706] = ~window[2][2];
assign temp[707] = ~window[2][3];
assign temp[708] = ~window[2][4];
assign temp[709] = window[2][5];
assign temp[710] = ~window[2][6];
assign temp[711] = window[2][7];
assign temp[712] = window[2][8];
assign temp[736] = window[3][0];
assign temp[737] = ~window[3][1];
assign temp[738] = ~window[3][2];
assign temp[739] = window[3][3];
assign temp[740] = window[3][4];
assign temp[741] = ~window[3][5];
assign temp[742] = window[3][6];
assign temp[743] = window[3][7];
assign temp[744] = ~window[3][8];
assign temp[768] = window[4][0];
assign temp[769] = ~window[4][1];
assign temp[770] = ~window[4][2];
assign temp[771] = ~window[4][3];
assign temp[772] = ~window[4][4];
assign temp[773] = ~window[4][5];
assign temp[774] = window[4][6];
assign temp[775] = ~window[4][7];
assign temp[776] = ~window[4][8];
assign temp[800] = ~window[5][0];
assign temp[801] = window[5][1];
assign temp[802] = ~window[5][2];
assign temp[803] = window[5][3];
assign temp[804] = window[5][4];
assign temp[805] = window[5][5];
assign temp[806] = ~window[5][6];
assign temp[807] = window[5][7];
assign temp[808] = window[5][8];
assign temp[832] = ~window[6][0];
assign temp[833] = window[6][1];
assign temp[834] = ~window[6][2];
assign temp[835] = ~window[6][3];
assign temp[836] = ~window[6][4];
assign temp[837] = window[6][5];
assign temp[838] = ~window[6][6];
assign temp[839] = ~window[6][7];
assign temp[840] = window[6][8];
assign temp[864] = window[7][0];
assign temp[865] = ~window[7][1];
assign temp[866] = ~window[7][2];
assign temp[867] = window[7][3];
assign temp[868] = ~window[7][4];
assign temp[869] = ~window[7][5];
assign temp[870] = window[7][6];
assign temp[871] = ~window[7][7];
assign temp[872] = ~window[7][8];
assign temp[896] = window[8][0];
assign temp[897] = ~window[8][1];
assign temp[898] = ~window[8][2];
assign temp[899] = ~window[8][3];
assign temp[900] = ~window[8][4];
assign temp[901] = window[8][5];
assign temp[902] = ~window[8][6];
assign temp[903] = ~window[8][7];
assign temp[904] = window[8][8];
assign temp[928] = window[9][0];
assign temp[929] = window[9][1];
assign temp[930] = ~window[9][2];
assign temp[931] = window[9][3];
assign temp[932] = ~window[9][4];
assign temp[933] = ~window[9][5];
assign temp[934] = window[9][6];
assign temp[935] = window[9][7];
assign temp[936] = window[9][8];
assign temp[960] = window[10][0];
assign temp[961] = window[10][1];
assign temp[962] = ~window[10][2];
assign temp[963] = window[10][3];
assign temp[964] = ~window[10][4];
assign temp[965] = ~window[10][5];
assign temp[966] = window[10][6];
assign temp[967] = ~window[10][7];
assign temp[968] = ~window[10][8];
assign temp[992] = window[11][0];
assign temp[993] = ~window[11][1];
assign temp[994] = window[11][2];
assign temp[995] = window[11][3];
assign temp[996] = ~window[11][4];
assign temp[997] = ~window[11][5];
assign temp[998] = window[11][6];
assign temp[999] = ~window[11][7];
assign temp[1000] = ~window[11][8];
assign temp[1024] = window[12][0];
assign temp[1025] = ~window[12][1];
assign temp[1026] = ~window[12][2];
assign temp[1027] = window[12][3];
assign temp[1028] = ~window[12][4];
assign temp[1029] = ~window[12][5];
assign temp[1030] = ~window[12][6];
assign temp[1031] = window[12][7];
assign temp[1032] = window[12][8];
assign temp[1056] = ~window[13][0];
assign temp[1057] = window[13][1];
assign temp[1058] = window[13][2];
assign temp[1059] = ~window[13][3];
assign temp[1060] = window[13][4];
assign temp[1061] = window[13][5];
assign temp[1062] = window[13][6];
assign temp[1063] = window[13][7];
assign temp[1064] = ~window[13][8];
assign temp[1088] = ~window[14][0];
assign temp[1089] = ~window[14][1];
assign temp[1090] = ~window[14][2];
assign temp[1091] = ~window[14][3];
assign temp[1092] = window[14][4];
assign temp[1093] = window[14][5];
assign temp[1094] = ~window[14][6];
assign temp[1095] = ~window[14][7];
assign temp[1096] = window[14][8];
assign temp[1120] = ~window[15][0];
assign temp[1121] = window[15][1];
assign temp[1122] = window[15][2];
assign temp[1123] = ~window[15][3];
assign temp[1124] = ~window[15][4];
assign temp[1125] = ~window[15][5];
assign temp[1126] = window[15][6];
assign temp[1127] = window[15][7];
assign temp[1128] = window[15][8];
assign temp[1152] = window[16][0];
assign temp[1153] = ~window[16][1];
assign temp[1154] = window[16][2];
assign temp[1155] = ~window[16][3];
assign temp[1156] = ~window[16][4];
assign temp[1157] = window[16][5];
assign temp[1158] = ~window[16][6];
assign temp[1159] = ~window[16][7];
assign temp[1160] = ~window[16][8];
assign temp[1184] = window[17][0];
assign temp[1185] = window[17][1];
assign temp[1186] = ~window[17][2];
assign temp[1187] = window[17][3];
assign temp[1188] = window[17][4];
assign temp[1189] = window[17][5];
assign temp[1190] = window[17][6];
assign temp[1191] = ~window[17][7];
assign temp[1192] = window[17][8];
assign temp[1216] = ~window[18][0];
assign temp[1217] = ~window[18][1];
assign temp[1218] = window[18][2];
assign temp[1219] = ~window[18][3];
assign temp[1220] = window[18][4];
assign temp[1221] = window[18][5];
assign temp[1222] = ~window[18][6];
assign temp[1223] = window[18][7];
assign temp[1224] = window[18][8];
assign temp[1248] = ~window[19][0];
assign temp[1249] = window[19][1];
assign temp[1250] = ~window[19][2];
assign temp[1251] = window[19][3];
assign temp[1252] = window[19][4];
assign temp[1253] = ~window[19][5];
assign temp[1254] = window[19][6];
assign temp[1255] = window[19][7];
assign temp[1256] = ~window[19][8];
assign temp[1280] = window[20][0];
assign temp[1281] = ~window[20][1];
assign temp[1282] = ~window[20][2];
assign temp[1283] = window[20][3];
assign temp[1284] = ~window[20][4];
assign temp[1285] = ~window[20][5];
assign temp[1286] = ~window[20][6];
assign temp[1287] = ~window[20][7];
assign temp[1288] = window[20][8];
assign temp[1312] = window[21][0];
assign temp[1313] = window[21][1];
assign temp[1314] = ~window[21][2];
assign temp[1315] = window[21][3];
assign temp[1316] = window[21][4];
assign temp[1317] = ~window[21][5];
assign temp[1318] = window[21][6];
assign temp[1319] = window[21][7];
assign temp[1320] = ~window[21][8];
assign temp[1344] = ~window[22][0];
assign temp[1345] = window[22][1];
assign temp[1346] = window[22][2];
assign temp[1347] = ~window[22][3];
assign temp[1348] = ~window[22][4];
assign temp[1349] = window[22][5];
assign temp[1350] = ~window[22][6];
assign temp[1351] = ~window[22][7];
assign temp[1352] = ~window[22][8];
assign temp[1376] = window[23][0];
assign temp[1377] = ~window[23][1];
assign temp[1378] = ~window[23][2];
assign temp[1379] = ~window[23][3];
assign temp[1380] = window[23][4];
assign temp[1381] = ~window[23][5];
assign temp[1382] = ~window[23][6];
assign temp[1383] = window[23][7];
assign temp[1384] = ~window[23][8];
assign temp[1408] = window[24][0];
assign temp[1409] = ~window[24][1];
assign temp[1410] = ~window[24][2];
assign temp[1411] = ~window[24][3];
assign temp[1412] = ~window[24][4];
assign temp[1413] = ~window[24][5];
assign temp[1414] = ~window[24][6];
assign temp[1415] = ~window[24][7];
assign temp[1416] = window[24][8];
assign temp[1440] = ~window[25][0];
assign temp[1441] = ~window[25][1];
assign temp[1442] = window[25][2];
assign temp[1443] = ~window[25][3];
assign temp[1444] = window[25][4];
assign temp[1445] = window[25][5];
assign temp[1446] = ~window[25][6];
assign temp[1447] = ~window[25][7];
assign temp[1448] = ~window[25][8];
assign temp[1472] = window[26][0];
assign temp[1473] = window[26][1];
assign temp[1474] = ~window[26][2];
assign temp[1475] = window[26][3];
assign temp[1476] = window[26][4];
assign temp[1477] = ~window[26][5];
assign temp[1478] = window[26][6];
assign temp[1479] = window[26][7];
assign temp[1480] = window[26][8];
assign temp[1504] = ~window[27][0];
assign temp[1505] = ~window[27][1];
assign temp[1506] = window[27][2];
assign temp[1507] = ~window[27][3];
assign temp[1508] = ~window[27][4];
assign temp[1509] = ~window[27][5];
assign temp[1510] = ~window[27][6];
assign temp[1511] = ~window[27][7];
assign temp[1512] = ~window[27][8];
assign temp[1536] = window[28][0];
assign temp[1537] = ~window[28][1];
assign temp[1538] = window[28][2];
assign temp[1539] = ~window[28][3];
assign temp[1540] = ~window[28][4];
assign temp[1541] = window[28][5];
assign temp[1542] = ~window[28][6];
assign temp[1543] = ~window[28][7];
assign temp[1544] = ~window[28][8];
assign temp[1568] = ~window[29][0];
assign temp[1569] = window[29][1];
assign temp[1570] = ~window[29][2];
assign temp[1571] = ~window[29][3];
assign temp[1572] = window[29][4];
assign temp[1573] = ~window[29][5];
assign temp[1574] = window[29][6];
assign temp[1575] = ~window[29][7];
assign temp[1576] = ~window[29][8];
assign temp[1600] = ~window[30][0];
assign temp[1601] = window[30][1];
assign temp[1602] = window[30][2];
assign temp[1603] = window[30][3];
assign temp[1604] = window[30][4];
assign temp[1605] = window[30][5];
assign temp[1606] = ~window[30][6];
assign temp[1607] = window[30][7];
assign temp[1608] = ~window[30][8];
assign temp[1632] = window[31][0];
assign temp[1633] = ~window[31][1];
assign temp[1634] = ~window[31][2];
assign temp[1635] = window[31][3];
assign temp[1636] = ~window[31][4];
assign temp[1637] = ~window[31][5];
assign temp[1638] = window[31][6];
assign temp[1639] = window[31][7];
assign temp[1640] = ~window[31][8];
assign temp[672] = ~window[0][0];
assign temp[673] = ~window[0][1];
assign temp[674] = ~window[0][2];
assign temp[675] = ~window[0][3];
assign temp[676] = window[0][4];
assign temp[677] = ~window[0][5];
assign temp[678] = ~window[0][6];
assign temp[679] = ~window[0][7];
assign temp[680] = ~window[0][8];
assign temp[704] = window[1][0];
assign temp[705] = ~window[1][1];
assign temp[706] = window[1][2];
assign temp[707] = ~window[1][3];
assign temp[708] = window[1][4];
assign temp[709] = window[1][5];
assign temp[710] = window[1][6];
assign temp[711] = window[1][7];
assign temp[712] = window[1][8];
assign temp[736] = window[2][0];
assign temp[737] = ~window[2][1];
assign temp[738] = ~window[2][2];
assign temp[739] = ~window[2][3];
assign temp[740] = ~window[2][4];
assign temp[741] = window[2][5];
assign temp[742] = ~window[2][6];
assign temp[743] = window[2][7];
assign temp[744] = ~window[2][8];
assign temp[768] = ~window[3][0];
assign temp[769] = ~window[3][1];
assign temp[770] = window[3][2];
assign temp[771] = ~window[3][3];
assign temp[772] = window[3][4];
assign temp[773] = window[3][5];
assign temp[774] = ~window[3][6];
assign temp[775] = window[3][7];
assign temp[776] = ~window[3][8];
assign temp[800] = ~window[4][0];
assign temp[801] = ~window[4][1];
assign temp[802] = ~window[4][2];
assign temp[803] = window[4][3];
assign temp[804] = ~window[4][4];
assign temp[805] = ~window[4][5];
assign temp[806] = ~window[4][6];
assign temp[807] = ~window[4][7];
assign temp[808] = ~window[4][8];
assign temp[832] = ~window[5][0];
assign temp[833] = window[5][1];
assign temp[834] = window[5][2];
assign temp[835] = ~window[5][3];
assign temp[836] = window[5][4];
assign temp[837] = ~window[5][5];
assign temp[838] = window[5][6];
assign temp[839] = window[5][7];
assign temp[840] = ~window[5][8];
assign temp[864] = window[6][0];
assign temp[865] = ~window[6][1];
assign temp[866] = ~window[6][2];
assign temp[867] = ~window[6][3];
assign temp[868] = ~window[6][4];
assign temp[869] = ~window[6][5];
assign temp[870] = ~window[6][6];
assign temp[871] = ~window[6][7];
assign temp[872] = window[6][8];
assign temp[896] = ~window[7][0];
assign temp[897] = window[7][1];
assign temp[898] = window[7][2];
assign temp[899] = ~window[7][3];
assign temp[900] = window[7][4];
assign temp[901] = window[7][5];
assign temp[902] = window[7][6];
assign temp[903] = ~window[7][7];
assign temp[904] = ~window[7][8];
assign temp[928] = ~window[8][0];
assign temp[929] = window[8][1];
assign temp[930] = window[8][2];
assign temp[931] = ~window[8][3];
assign temp[932] = ~window[8][4];
assign temp[933] = ~window[8][5];
assign temp[934] = ~window[8][6];
assign temp[935] = ~window[8][7];
assign temp[936] = ~window[8][8];
assign temp[960] = ~window[9][0];
assign temp[961] = ~window[9][1];
assign temp[962] = window[9][2];
assign temp[963] = ~window[9][3];
assign temp[964] = window[9][4];
assign temp[965] = window[9][5];
assign temp[966] = ~window[9][6];
assign temp[967] = window[9][7];
assign temp[968] = ~window[9][8];
assign temp[992] = ~window[10][0];
assign temp[993] = window[10][1];
assign temp[994] = ~window[10][2];
assign temp[995] = ~window[10][3];
assign temp[996] = window[10][4];
assign temp[997] = window[10][5];
assign temp[998] = ~window[10][6];
assign temp[999] = window[10][7];
assign temp[1000] = ~window[10][8];
assign temp[1024] = ~window[11][0];
assign temp[1025] = window[11][1];
assign temp[1026] = ~window[11][2];
assign temp[1027] = ~window[11][3];
assign temp[1028] = window[11][4];
assign temp[1029] = window[11][5];
assign temp[1030] = window[11][6];
assign temp[1031] = window[11][7];
assign temp[1032] = window[11][8];
assign temp[1056] = window[12][0];
assign temp[1057] = window[12][1];
assign temp[1058] = ~window[12][2];
assign temp[1059] = ~window[12][3];
assign temp[1060] = ~window[12][4];
assign temp[1061] = ~window[12][5];
assign temp[1062] = ~window[12][6];
assign temp[1063] = window[12][7];
assign temp[1064] = window[12][8];
assign temp[1088] = ~window[13][0];
assign temp[1089] = window[13][1];
assign temp[1090] = window[13][2];
assign temp[1091] = window[13][3];
assign temp[1092] = window[13][4];
assign temp[1093] = window[13][5];
assign temp[1094] = window[13][6];
assign temp[1095] = window[13][7];
assign temp[1096] = window[13][8];
assign temp[1120] = ~window[14][0];
assign temp[1121] = ~window[14][1];
assign temp[1122] = window[14][2];
assign temp[1123] = ~window[14][3];
assign temp[1124] = ~window[14][4];
assign temp[1125] = ~window[14][5];
assign temp[1126] = window[14][6];
assign temp[1127] = ~window[14][7];
assign temp[1128] = ~window[14][8];
assign temp[1152] = window[15][0];
assign temp[1153] = window[15][1];
assign temp[1154] = ~window[15][2];
assign temp[1155] = window[15][3];
assign temp[1156] = ~window[15][4];
assign temp[1157] = ~window[15][5];
assign temp[1158] = ~window[15][6];
assign temp[1159] = ~window[15][7];
assign temp[1160] = window[15][8];
assign temp[1184] = window[16][0];
assign temp[1185] = window[16][1];
assign temp[1186] = ~window[16][2];
assign temp[1187] = window[16][3];
assign temp[1188] = window[16][4];
assign temp[1189] = ~window[16][5];
assign temp[1190] = window[16][6];
assign temp[1191] = window[16][7];
assign temp[1192] = ~window[16][8];
assign temp[1216] = window[17][0];
assign temp[1217] = window[17][1];
assign temp[1218] = window[17][2];
assign temp[1219] = ~window[17][3];
assign temp[1220] = window[17][4];
assign temp[1221] = window[17][5];
assign temp[1222] = window[17][6];
assign temp[1223] = window[17][7];
assign temp[1224] = window[17][8];
assign temp[1248] = ~window[18][0];
assign temp[1249] = ~window[18][1];
assign temp[1250] = ~window[18][2];
assign temp[1251] = ~window[18][3];
assign temp[1252] = ~window[18][4];
assign temp[1253] = window[18][5];
assign temp[1254] = ~window[18][6];
assign temp[1255] = window[18][7];
assign temp[1256] = ~window[18][8];
assign temp[1280] = ~window[19][0];
assign temp[1281] = ~window[19][1];
assign temp[1282] = ~window[19][2];
assign temp[1283] = ~window[19][3];
assign temp[1284] = window[19][4];
assign temp[1285] = window[19][5];
assign temp[1286] = window[19][6];
assign temp[1287] = window[19][7];
assign temp[1288] = window[19][8];
assign temp[1312] = ~window[20][0];
assign temp[1313] = ~window[20][1];
assign temp[1314] = window[20][2];
assign temp[1315] = ~window[20][3];
assign temp[1316] = window[20][4];
assign temp[1317] = window[20][5];
assign temp[1318] = window[20][6];
assign temp[1319] = window[20][7];
assign temp[1320] = ~window[20][8];
assign temp[1344] = ~window[21][0];
assign temp[1345] = ~window[21][1];
assign temp[1346] = ~window[21][2];
assign temp[1347] = ~window[21][3];
assign temp[1348] = window[21][4];
assign temp[1349] = window[21][5];
assign temp[1350] = window[21][6];
assign temp[1351] = window[21][7];
assign temp[1352] = ~window[21][8];
assign temp[1376] = window[22][0];
assign temp[1377] = window[22][1];
assign temp[1378] = ~window[22][2];
assign temp[1379] = window[22][3];
assign temp[1380] = ~window[22][4];
assign temp[1381] = ~window[22][5];
assign temp[1382] = ~window[22][6];
assign temp[1383] = ~window[22][7];
assign temp[1384] = ~window[22][8];
assign temp[1408] = window[23][0];
assign temp[1409] = ~window[23][1];
assign temp[1410] = window[23][2];
assign temp[1411] = ~window[23][3];
assign temp[1412] = window[23][4];
assign temp[1413] = ~window[23][5];
assign temp[1414] = window[23][6];
assign temp[1415] = window[23][7];
assign temp[1416] = ~window[23][8];
assign temp[1440] = window[24][0];
assign temp[1441] = ~window[24][1];
assign temp[1442] = window[24][2];
assign temp[1443] = ~window[24][3];
assign temp[1444] = ~window[24][4];
assign temp[1445] = window[24][5];
assign temp[1446] = ~window[24][6];
assign temp[1447] = window[24][7];
assign temp[1448] = ~window[24][8];
assign temp[1472] = window[25][0];
assign temp[1473] = window[25][1];
assign temp[1474] = window[25][2];
assign temp[1475] = window[25][3];
assign temp[1476] = window[25][4];
assign temp[1477] = ~window[25][5];
assign temp[1478] = window[25][6];
assign temp[1479] = ~window[25][7];
assign temp[1480] = ~window[25][8];
assign temp[1504] = ~window[26][0];
assign temp[1505] = window[26][1];
assign temp[1506] = ~window[26][2];
assign temp[1507] = ~window[26][3];
assign temp[1508] = ~window[26][4];
assign temp[1509] = window[26][5];
assign temp[1510] = ~window[26][6];
assign temp[1511] = window[26][7];
assign temp[1512] = window[26][8];
assign temp[1536] = ~window[27][0];
assign temp[1537] = ~window[27][1];
assign temp[1538] = ~window[27][2];
assign temp[1539] = window[27][3];
assign temp[1540] = window[27][4];
assign temp[1541] = ~window[27][5];
assign temp[1542] = window[27][6];
assign temp[1543] = ~window[27][7];
assign temp[1544] = ~window[27][8];
assign temp[1568] = window[28][0];
assign temp[1569] = window[28][1];
assign temp[1570] = window[28][2];
assign temp[1571] = window[28][3];
assign temp[1572] = window[28][4];
assign temp[1573] = ~window[28][5];
assign temp[1574] = ~window[28][6];
assign temp[1575] = window[28][7];
assign temp[1576] = ~window[28][8];
assign temp[1600] = ~window[29][0];
assign temp[1601] = window[29][1];
assign temp[1602] = window[29][2];
assign temp[1603] = window[29][3];
assign temp[1604] = window[29][4];
assign temp[1605] = window[29][5];
assign temp[1606] = window[29][6];
assign temp[1607] = window[29][7];
assign temp[1608] = ~window[29][8];
assign temp[1632] = window[30][0];
assign temp[1633] = window[30][1];
assign temp[1634] = window[30][2];
assign temp[1635] = window[30][3];
assign temp[1636] = window[30][4];
assign temp[1637] = window[30][5];
assign temp[1638] = window[30][6];
assign temp[1639] = window[30][7];
assign temp[1640] = ~window[30][8];
assign temp[1664] = window[31][0];
assign temp[1665] = window[31][1];
assign temp[1666] = ~window[31][2];
assign temp[1667] = ~window[31][3];
assign temp[1668] = ~window[31][4];
assign temp[1669] = window[31][5];
assign temp[1670] = ~window[31][6];
assign temp[1671] = window[31][7];
assign temp[1672] = ~window[31][8];
assign temp[704] = ~window[0][0];
assign temp[705] = ~window[0][1];
assign temp[706] = ~window[0][2];
assign temp[707] = ~window[0][3];
assign temp[708] = ~window[0][4];
assign temp[709] = ~window[0][5];
assign temp[710] = window[0][6];
assign temp[711] = window[0][7];
assign temp[712] = window[0][8];
assign temp[736] = ~window[1][0];
assign temp[737] = ~window[1][1];
assign temp[738] = ~window[1][2];
assign temp[739] = window[1][3];
assign temp[740] = ~window[1][4];
assign temp[741] = ~window[1][5];
assign temp[742] = window[1][6];
assign temp[743] = window[1][7];
assign temp[744] = ~window[1][8];
assign temp[768] = ~window[2][0];
assign temp[769] = ~window[2][1];
assign temp[770] = window[2][2];
assign temp[771] = ~window[2][3];
assign temp[772] = ~window[2][4];
assign temp[773] = ~window[2][5];
assign temp[774] = window[2][6];
assign temp[775] = window[2][7];
assign temp[776] = ~window[2][8];
assign temp[800] = ~window[3][0];
assign temp[801] = ~window[3][1];
assign temp[802] = ~window[3][2];
assign temp[803] = ~window[3][3];
assign temp[804] = ~window[3][4];
assign temp[805] = ~window[3][5];
assign temp[806] = window[3][6];
assign temp[807] = window[3][7];
assign temp[808] = window[3][8];
assign temp[832] = ~window[4][0];
assign temp[833] = ~window[4][1];
assign temp[834] = window[4][2];
assign temp[835] = ~window[4][3];
assign temp[836] = window[4][4];
assign temp[837] = window[4][5];
assign temp[838] = window[4][6];
assign temp[839] = window[4][7];
assign temp[840] = window[4][8];
assign temp[864] = ~window[5][0];
assign temp[865] = ~window[5][1];
assign temp[866] = ~window[5][2];
assign temp[867] = window[5][3];
assign temp[868] = ~window[5][4];
assign temp[869] = window[5][5];
assign temp[870] = window[5][6];
assign temp[871] = window[5][7];
assign temp[872] = window[5][8];
assign temp[896] = ~window[6][0];
assign temp[897] = ~window[6][1];
assign temp[898] = window[6][2];
assign temp[899] = ~window[6][3];
assign temp[900] = window[6][4];
assign temp[901] = window[6][5];
assign temp[902] = window[6][6];
assign temp[903] = ~window[6][7];
assign temp[904] = ~window[6][8];
assign temp[928] = window[7][0];
assign temp[929] = ~window[7][1];
assign temp[930] = ~window[7][2];
assign temp[931] = window[7][3];
assign temp[932] = window[7][4];
assign temp[933] = window[7][5];
assign temp[934] = window[7][6];
assign temp[935] = window[7][7];
assign temp[936] = window[7][8];
assign temp[960] = ~window[8][0];
assign temp[961] = ~window[8][1];
assign temp[962] = ~window[8][2];
assign temp[963] = ~window[8][3];
assign temp[964] = window[8][4];
assign temp[965] = window[8][5];
assign temp[966] = window[8][6];
assign temp[967] = window[8][7];
assign temp[968] = window[8][8];
assign temp[992] = ~window[9][0];
assign temp[993] = ~window[9][1];
assign temp[994] = ~window[9][2];
assign temp[995] = window[9][3];
assign temp[996] = window[9][4];
assign temp[997] = ~window[9][5];
assign temp[998] = window[9][6];
assign temp[999] = window[9][7];
assign temp[1000] = window[9][8];
assign temp[1024] = window[10][0];
assign temp[1025] = window[10][1];
assign temp[1026] = ~window[10][2];
assign temp[1027] = window[10][3];
assign temp[1028] = window[10][4];
assign temp[1029] = window[10][5];
assign temp[1030] = window[10][6];
assign temp[1031] = window[10][7];
assign temp[1032] = window[10][8];
assign temp[1056] = ~window[11][0];
assign temp[1057] = ~window[11][1];
assign temp[1058] = window[11][2];
assign temp[1059] = ~window[11][3];
assign temp[1060] = window[11][4];
assign temp[1061] = window[11][5];
assign temp[1062] = window[11][6];
assign temp[1063] = ~window[11][7];
assign temp[1064] = window[11][8];
assign temp[1088] = ~window[12][0];
assign temp[1089] = window[12][1];
assign temp[1090] = window[12][2];
assign temp[1091] = ~window[12][3];
assign temp[1092] = ~window[12][4];
assign temp[1093] = window[12][5];
assign temp[1094] = window[12][6];
assign temp[1095] = window[12][7];
assign temp[1096] = ~window[12][8];
assign temp[1120] = ~window[13][0];
assign temp[1121] = window[13][1];
assign temp[1122] = window[13][2];
assign temp[1123] = ~window[13][3];
assign temp[1124] = window[13][4];
assign temp[1125] = window[13][5];
assign temp[1126] = ~window[13][6];
assign temp[1127] = window[13][7];
assign temp[1128] = ~window[13][8];
assign temp[1152] = ~window[14][0];
assign temp[1153] = ~window[14][1];
assign temp[1154] = ~window[14][2];
assign temp[1155] = ~window[14][3];
assign temp[1156] = ~window[14][4];
assign temp[1157] = window[14][5];
assign temp[1158] = window[14][6];
assign temp[1159] = window[14][7];
assign temp[1160] = window[14][8];
assign temp[1184] = window[15][0];
assign temp[1185] = ~window[15][1];
assign temp[1186] = window[15][2];
assign temp[1187] = window[15][3];
assign temp[1188] = ~window[15][4];
assign temp[1189] = window[15][5];
assign temp[1190] = window[15][6];
assign temp[1191] = ~window[15][7];
assign temp[1192] = ~window[15][8];
assign temp[1216] = window[16][0];
assign temp[1217] = ~window[16][1];
assign temp[1218] = ~window[16][2];
assign temp[1219] = ~window[16][3];
assign temp[1220] = window[16][4];
assign temp[1221] = window[16][5];
assign temp[1222] = ~window[16][6];
assign temp[1223] = window[16][7];
assign temp[1224] = window[16][8];
assign temp[1248] = ~window[17][0];
assign temp[1249] = ~window[17][1];
assign temp[1250] = ~window[17][2];
assign temp[1251] = window[17][3];
assign temp[1252] = ~window[17][4];
assign temp[1253] = ~window[17][5];
assign temp[1254] = window[17][6];
assign temp[1255] = window[17][7];
assign temp[1256] = window[17][8];
assign temp[1280] = window[18][0];
assign temp[1281] = ~window[18][1];
assign temp[1282] = window[18][2];
assign temp[1283] = ~window[18][3];
assign temp[1284] = window[18][4];
assign temp[1285] = ~window[18][5];
assign temp[1286] = ~window[18][6];
assign temp[1287] = ~window[18][7];
assign temp[1288] = ~window[18][8];
assign temp[1312] = window[19][0];
assign temp[1313] = window[19][1];
assign temp[1314] = window[19][2];
assign temp[1315] = ~window[19][3];
assign temp[1316] = ~window[19][4];
assign temp[1317] = ~window[19][5];
assign temp[1318] = ~window[19][6];
assign temp[1319] = ~window[19][7];
assign temp[1320] = ~window[19][8];
assign temp[1344] = ~window[20][0];
assign temp[1345] = ~window[20][1];
assign temp[1346] = ~window[20][2];
assign temp[1347] = ~window[20][3];
assign temp[1348] = ~window[20][4];
assign temp[1349] = ~window[20][5];
assign temp[1350] = window[20][6];
assign temp[1351] = window[20][7];
assign temp[1352] = window[20][8];
assign temp[1376] = window[21][0];
assign temp[1377] = window[21][1];
assign temp[1378] = window[21][2];
assign temp[1379] = window[21][3];
assign temp[1380] = ~window[21][4];
assign temp[1381] = window[21][5];
assign temp[1382] = window[21][6];
assign temp[1383] = ~window[21][7];
assign temp[1384] = window[21][8];
assign temp[1408] = window[22][0];
assign temp[1409] = window[22][1];
assign temp[1410] = window[22][2];
assign temp[1411] = ~window[22][3];
assign temp[1412] = window[22][4];
assign temp[1413] = window[22][5];
assign temp[1414] = ~window[22][6];
assign temp[1415] = ~window[22][7];
assign temp[1416] = ~window[22][8];
assign temp[1440] = ~window[23][0];
assign temp[1441] = ~window[23][1];
assign temp[1442] = ~window[23][2];
assign temp[1443] = window[23][3];
assign temp[1444] = ~window[23][4];
assign temp[1445] = ~window[23][5];
assign temp[1446] = window[23][6];
assign temp[1447] = ~window[23][7];
assign temp[1448] = window[23][8];
assign temp[1472] = ~window[24][0];
assign temp[1473] = ~window[24][1];
assign temp[1474] = ~window[24][2];
assign temp[1475] = ~window[24][3];
assign temp[1476] = ~window[24][4];
assign temp[1477] = ~window[24][5];
assign temp[1478] = window[24][6];
assign temp[1479] = window[24][7];
assign temp[1480] = window[24][8];
assign temp[1504] = ~window[25][0];
assign temp[1505] = ~window[25][1];
assign temp[1506] = ~window[25][2];
assign temp[1507] = ~window[25][3];
assign temp[1508] = window[25][4];
assign temp[1509] = ~window[25][5];
assign temp[1510] = window[25][6];
assign temp[1511] = window[25][7];
assign temp[1512] = window[25][8];
assign temp[1536] = ~window[26][0];
assign temp[1537] = window[26][1];
assign temp[1538] = window[26][2];
assign temp[1539] = window[26][3];
assign temp[1540] = ~window[26][4];
assign temp[1541] = ~window[26][5];
assign temp[1542] = window[26][6];
assign temp[1543] = ~window[26][7];
assign temp[1544] = window[26][8];
assign temp[1568] = window[27][0];
assign temp[1569] = window[27][1];
assign temp[1570] = ~window[27][2];
assign temp[1571] = window[27][3];
assign temp[1572] = window[27][4];
assign temp[1573] = window[27][5];
assign temp[1574] = ~window[27][6];
assign temp[1575] = window[27][7];
assign temp[1576] = window[27][8];
assign temp[1600] = window[28][0];
assign temp[1601] = window[28][1];
assign temp[1602] = window[28][2];
assign temp[1603] = ~window[28][3];
assign temp[1604] = ~window[28][4];
assign temp[1605] = window[28][5];
assign temp[1606] = window[28][6];
assign temp[1607] = window[28][7];
assign temp[1608] = window[28][8];
assign temp[1632] = window[29][0];
assign temp[1633] = window[29][1];
assign temp[1634] = ~window[29][2];
assign temp[1635] = ~window[29][3];
assign temp[1636] = ~window[29][4];
assign temp[1637] = window[29][5];
assign temp[1638] = ~window[29][6];
assign temp[1639] = ~window[29][7];
assign temp[1640] = window[29][8];
assign temp[1664] = ~window[30][0];
assign temp[1665] = ~window[30][1];
assign temp[1666] = window[30][2];
assign temp[1667] = ~window[30][3];
assign temp[1668] = ~window[30][4];
assign temp[1669] = ~window[30][5];
assign temp[1670] = ~window[30][6];
assign temp[1671] = ~window[30][7];
assign temp[1672] = ~window[30][8];
assign temp[1696] = ~window[31][0];
assign temp[1697] = ~window[31][1];
assign temp[1698] = ~window[31][2];
assign temp[1699] = window[31][3];
assign temp[1700] = ~window[31][4];
assign temp[1701] = window[31][5];
assign temp[1702] = window[31][6];
assign temp[1703] = window[31][7];
assign temp[1704] = window[31][8];
assign temp[736] = ~window[0][0];
assign temp[737] = window[0][1];
assign temp[738] = ~window[0][2];
assign temp[739] = window[0][3];
assign temp[740] = window[0][4];
assign temp[741] = ~window[0][5];
assign temp[742] = window[0][6];
assign temp[743] = window[0][7];
assign temp[744] = ~window[0][8];
assign temp[768] = ~window[1][0];
assign temp[769] = window[1][1];
assign temp[770] = ~window[1][2];
assign temp[771] = window[1][3];
assign temp[772] = window[1][4];
assign temp[773] = window[1][5];
assign temp[774] = ~window[1][6];
assign temp[775] = ~window[1][7];
assign temp[776] = ~window[1][8];
assign temp[800] = window[2][0];
assign temp[801] = ~window[2][1];
assign temp[802] = window[2][2];
assign temp[803] = window[2][3];
assign temp[804] = window[2][4];
assign temp[805] = window[2][5];
assign temp[806] = window[2][6];
assign temp[807] = window[2][7];
assign temp[808] = ~window[2][8];
assign temp[832] = ~window[3][0];
assign temp[833] = ~window[3][1];
assign temp[834] = window[3][2];
assign temp[835] = ~window[3][3];
assign temp[836] = ~window[3][4];
assign temp[837] = window[3][5];
assign temp[838] = ~window[3][6];
assign temp[839] = ~window[3][7];
assign temp[840] = ~window[3][8];
assign temp[864] = ~window[4][0];
assign temp[865] = ~window[4][1];
assign temp[866] = ~window[4][2];
assign temp[867] = window[4][3];
assign temp[868] = window[4][4];
assign temp[869] = ~window[4][5];
assign temp[870] = window[4][6];
assign temp[871] = window[4][7];
assign temp[872] = window[4][8];
assign temp[896] = ~window[5][0];
assign temp[897] = window[5][1];
assign temp[898] = window[5][2];
assign temp[899] = window[5][3];
assign temp[900] = ~window[5][4];
assign temp[901] = ~window[5][5];
assign temp[902] = ~window[5][6];
assign temp[903] = ~window[5][7];
assign temp[904] = ~window[5][8];
assign temp[928] = window[6][0];
assign temp[929] = ~window[6][1];
assign temp[930] = ~window[6][2];
assign temp[931] = window[6][3];
assign temp[932] = window[6][4];
assign temp[933] = window[6][5];
assign temp[934] = window[6][6];
assign temp[935] = window[6][7];
assign temp[936] = window[6][8];
assign temp[960] = ~window[7][0];
assign temp[961] = window[7][1];
assign temp[962] = window[7][2];
assign temp[963] = ~window[7][3];
assign temp[964] = window[7][4];
assign temp[965] = ~window[7][5];
assign temp[966] = window[7][6];
assign temp[967] = window[7][7];
assign temp[968] = ~window[7][8];
assign temp[992] = ~window[8][0];
assign temp[993] = window[8][1];
assign temp[994] = window[8][2];
assign temp[995] = window[8][3];
assign temp[996] = window[8][4];
assign temp[997] = window[8][5];
assign temp[998] = window[8][6];
assign temp[999] = window[8][7];
assign temp[1000] = ~window[8][8];
assign temp[1024] = ~window[9][0];
assign temp[1025] = window[9][1];
assign temp[1026] = ~window[9][2];
assign temp[1027] = ~window[9][3];
assign temp[1028] = window[9][4];
assign temp[1029] = window[9][5];
assign temp[1030] = ~window[9][6];
assign temp[1031] = ~window[9][7];
assign temp[1032] = ~window[9][8];
assign temp[1056] = ~window[10][0];
assign temp[1057] = ~window[10][1];
assign temp[1058] = ~window[10][2];
assign temp[1059] = ~window[10][3];
assign temp[1060] = ~window[10][4];
assign temp[1061] = ~window[10][5];
assign temp[1062] = window[10][6];
assign temp[1063] = window[10][7];
assign temp[1064] = ~window[10][8];
assign temp[1088] = ~window[11][0];
assign temp[1089] = ~window[11][1];
assign temp[1090] = ~window[11][2];
assign temp[1091] = ~window[11][3];
assign temp[1092] = ~window[11][4];
assign temp[1093] = ~window[11][5];
assign temp[1094] = window[11][6];
assign temp[1095] = window[11][7];
assign temp[1096] = window[11][8];
assign temp[1120] = ~window[12][0];
assign temp[1121] = ~window[12][1];
assign temp[1122] = ~window[12][2];
assign temp[1123] = window[12][3];
assign temp[1124] = window[12][4];
assign temp[1125] = ~window[12][5];
assign temp[1126] = ~window[12][6];
assign temp[1127] = window[12][7];
assign temp[1128] = window[12][8];
assign temp[1152] = ~window[13][0];
assign temp[1153] = window[13][1];
assign temp[1154] = window[13][2];
assign temp[1155] = ~window[13][3];
assign temp[1156] = ~window[13][4];
assign temp[1157] = ~window[13][5];
assign temp[1158] = ~window[13][6];
assign temp[1159] = ~window[13][7];
assign temp[1160] = ~window[13][8];
assign temp[1184] = ~window[14][0];
assign temp[1185] = ~window[14][1];
assign temp[1186] = ~window[14][2];
assign temp[1187] = window[14][3];
assign temp[1188] = window[14][4];
assign temp[1189] = ~window[14][5];
assign temp[1190] = ~window[14][6];
assign temp[1191] = window[14][7];
assign temp[1192] = ~window[14][8];
assign temp[1216] = window[15][0];
assign temp[1217] = ~window[15][1];
assign temp[1218] = ~window[15][2];
assign temp[1219] = window[15][3];
assign temp[1220] = ~window[15][4];
assign temp[1221] = ~window[15][5];
assign temp[1222] = window[15][6];
assign temp[1223] = window[15][7];
assign temp[1224] = window[15][8];
assign temp[1248] = window[16][0];
assign temp[1249] = window[16][1];
assign temp[1250] = window[16][2];
assign temp[1251] = ~window[16][3];
assign temp[1252] = ~window[16][4];
assign temp[1253] = ~window[16][5];
assign temp[1254] = window[16][6];
assign temp[1255] = window[16][7];
assign temp[1256] = ~window[16][8];
assign temp[1280] = ~window[17][0];
assign temp[1281] = ~window[17][1];
assign temp[1282] = window[17][2];
assign temp[1283] = ~window[17][3];
assign temp[1284] = window[17][4];
assign temp[1285] = window[17][5];
assign temp[1286] = ~window[17][6];
assign temp[1287] = window[17][7];
assign temp[1288] = ~window[17][8];
assign temp[1312] = window[18][0];
assign temp[1313] = window[18][1];
assign temp[1314] = ~window[18][2];
assign temp[1315] = window[18][3];
assign temp[1316] = window[18][4];
assign temp[1317] = window[18][5];
assign temp[1318] = ~window[18][6];
assign temp[1319] = ~window[18][7];
assign temp[1320] = ~window[18][8];
assign temp[1344] = window[19][0];
assign temp[1345] = window[19][1];
assign temp[1346] = ~window[19][2];
assign temp[1347] = ~window[19][3];
assign temp[1348] = ~window[19][4];
assign temp[1349] = window[19][5];
assign temp[1350] = ~window[19][6];
assign temp[1351] = ~window[19][7];
assign temp[1352] = window[19][8];
assign temp[1376] = window[20][0];
assign temp[1377] = ~window[20][1];
assign temp[1378] = window[20][2];
assign temp[1379] = ~window[20][3];
assign temp[1380] = window[20][4];
assign temp[1381] = ~window[20][5];
assign temp[1382] = ~window[20][6];
assign temp[1383] = ~window[20][7];
assign temp[1384] = ~window[20][8];
assign temp[1408] = ~window[21][0];
assign temp[1409] = window[21][1];
assign temp[1410] = window[21][2];
assign temp[1411] = ~window[21][3];
assign temp[1412] = ~window[21][4];
assign temp[1413] = ~window[21][5];
assign temp[1414] = ~window[21][6];
assign temp[1415] = window[21][7];
assign temp[1416] = ~window[21][8];
assign temp[1440] = ~window[22][0];
assign temp[1441] = ~window[22][1];
assign temp[1442] = ~window[22][2];
assign temp[1443] = ~window[22][3];
assign temp[1444] = window[22][4];
assign temp[1445] = window[22][5];
assign temp[1446] = window[22][6];
assign temp[1447] = window[22][7];
assign temp[1448] = window[22][8];
assign temp[1472] = ~window[23][0];
assign temp[1473] = window[23][1];
assign temp[1474] = ~window[23][2];
assign temp[1475] = ~window[23][3];
assign temp[1476] = ~window[23][4];
assign temp[1477] = ~window[23][5];
assign temp[1478] = ~window[23][6];
assign temp[1479] = ~window[23][7];
assign temp[1480] = ~window[23][8];
assign temp[1504] = window[24][0];
assign temp[1505] = ~window[24][1];
assign temp[1506] = ~window[24][2];
assign temp[1507] = window[24][3];
assign temp[1508] = window[24][4];
assign temp[1509] = window[24][5];
assign temp[1510] = ~window[24][6];
assign temp[1511] = window[24][7];
assign temp[1512] = window[24][8];
assign temp[1536] = window[25][0];
assign temp[1537] = ~window[25][1];
assign temp[1538] = ~window[25][2];
assign temp[1539] = ~window[25][3];
assign temp[1540] = window[25][4];
assign temp[1541] = ~window[25][5];
assign temp[1542] = ~window[25][6];
assign temp[1543] = ~window[25][7];
assign temp[1544] = ~window[25][8];
assign temp[1568] = ~window[26][0];
assign temp[1569] = ~window[26][1];
assign temp[1570] = ~window[26][2];
assign temp[1571] = window[26][3];
assign temp[1572] = window[26][4];
assign temp[1573] = ~window[26][5];
assign temp[1574] = ~window[26][6];
assign temp[1575] = window[26][7];
assign temp[1576] = window[26][8];
assign temp[1600] = ~window[27][0];
assign temp[1601] = window[27][1];
assign temp[1602] = window[27][2];
assign temp[1603] = ~window[27][3];
assign temp[1604] = ~window[27][4];
assign temp[1605] = ~window[27][5];
assign temp[1606] = window[27][6];
assign temp[1607] = window[27][7];
assign temp[1608] = window[27][8];
assign temp[1632] = ~window[28][0];
assign temp[1633] = window[28][1];
assign temp[1634] = ~window[28][2];
assign temp[1635] = ~window[28][3];
assign temp[1636] = ~window[28][4];
assign temp[1637] = ~window[28][5];
assign temp[1638] = ~window[28][6];
assign temp[1639] = ~window[28][7];
assign temp[1640] = ~window[28][8];
assign temp[1664] = ~window[29][0];
assign temp[1665] = ~window[29][1];
assign temp[1666] = ~window[29][2];
assign temp[1667] = ~window[29][3];
assign temp[1668] = window[29][4];
assign temp[1669] = ~window[29][5];
assign temp[1670] = window[29][6];
assign temp[1671] = window[29][7];
assign temp[1672] = window[29][8];
assign temp[1696] = ~window[30][0];
assign temp[1697] = window[30][1];
assign temp[1698] = ~window[30][2];
assign temp[1699] = ~window[30][3];
assign temp[1700] = ~window[30][4];
assign temp[1701] = ~window[30][5];
assign temp[1702] = ~window[30][6];
assign temp[1703] = ~window[30][7];
assign temp[1704] = ~window[30][8];
assign temp[1728] = ~window[31][0];
assign temp[1729] = ~window[31][1];
assign temp[1730] = ~window[31][2];
assign temp[1731] = window[31][3];
assign temp[1732] = window[31][4];
assign temp[1733] = window[31][5];
assign temp[1734] = window[31][6];
assign temp[1735] = ~window[31][7];
assign temp[1736] = ~window[31][8];
assign temp[768] = ~window[0][0];
assign temp[769] = ~window[0][1];
assign temp[770] = ~window[0][2];
assign temp[771] = window[0][3];
assign temp[772] = ~window[0][4];
assign temp[773] = ~window[0][5];
assign temp[774] = window[0][6];
assign temp[775] = window[0][7];
assign temp[776] = window[0][8];
assign temp[800] = window[1][0];
assign temp[801] = ~window[1][1];
assign temp[802] = ~window[1][2];
assign temp[803] = window[1][3];
assign temp[804] = window[1][4];
assign temp[805] = window[1][5];
assign temp[806] = window[1][6];
assign temp[807] = window[1][7];
assign temp[808] = ~window[1][8];
assign temp[832] = ~window[2][0];
assign temp[833] = ~window[2][1];
assign temp[834] = ~window[2][2];
assign temp[835] = ~window[2][3];
assign temp[836] = ~window[2][4];
assign temp[837] = window[2][5];
assign temp[838] = ~window[2][6];
assign temp[839] = window[2][7];
assign temp[840] = window[2][8];
assign temp[864] = window[3][0];
assign temp[865] = ~window[3][1];
assign temp[866] = ~window[3][2];
assign temp[867] = window[3][3];
assign temp[868] = ~window[3][4];
assign temp[869] = window[3][5];
assign temp[870] = window[3][6];
assign temp[871] = window[3][7];
assign temp[872] = window[3][8];
assign temp[896] = window[4][0];
assign temp[897] = window[4][1];
assign temp[898] = window[4][2];
assign temp[899] = window[4][3];
assign temp[900] = window[4][4];
assign temp[901] = ~window[4][5];
assign temp[902] = window[4][6];
assign temp[903] = window[4][7];
assign temp[904] = ~window[4][8];
assign temp[928] = ~window[5][0];
assign temp[929] = ~window[5][1];
assign temp[930] = ~window[5][2];
assign temp[931] = window[5][3];
assign temp[932] = ~window[5][4];
assign temp[933] = ~window[5][5];
assign temp[934] = window[5][6];
assign temp[935] = ~window[5][7];
assign temp[936] = window[5][8];
assign temp[960] = window[6][0];
assign temp[961] = window[6][1];
assign temp[962] = window[6][2];
assign temp[963] = ~window[6][3];
assign temp[964] = ~window[6][4];
assign temp[965] = ~window[6][5];
assign temp[966] = window[6][6];
assign temp[967] = window[6][7];
assign temp[968] = window[6][8];
assign temp[992] = window[7][0];
assign temp[993] = window[7][1];
assign temp[994] = window[7][2];
assign temp[995] = window[7][3];
assign temp[996] = window[7][4];
assign temp[997] = window[7][5];
assign temp[998] = window[7][6];
assign temp[999] = ~window[7][7];
assign temp[1000] = ~window[7][8];
assign temp[1024] = ~window[8][0];
assign temp[1025] = ~window[8][1];
assign temp[1026] = ~window[8][2];
assign temp[1027] = window[8][3];
assign temp[1028] = ~window[8][4];
assign temp[1029] = window[8][5];
assign temp[1030] = ~window[8][6];
assign temp[1031] = window[8][7];
assign temp[1032] = window[8][8];
assign temp[1056] = window[9][0];
assign temp[1057] = ~window[9][1];
assign temp[1058] = ~window[9][2];
assign temp[1059] = window[9][3];
assign temp[1060] = window[9][4];
assign temp[1061] = window[9][5];
assign temp[1062] = window[9][6];
assign temp[1063] = window[9][7];
assign temp[1064] = window[9][8];
assign temp[1088] = window[10][0];
assign temp[1089] = ~window[10][1];
assign temp[1090] = ~window[10][2];
assign temp[1091] = window[10][3];
assign temp[1092] = window[10][4];
assign temp[1093] = window[10][5];
assign temp[1094] = window[10][6];
assign temp[1095] = ~window[10][7];
assign temp[1096] = ~window[10][8];
assign temp[1120] = ~window[11][0];
assign temp[1121] = window[11][1];
assign temp[1122] = window[11][2];
assign temp[1123] = ~window[11][3];
assign temp[1124] = ~window[11][4];
assign temp[1125] = window[11][5];
assign temp[1126] = window[11][6];
assign temp[1127] = ~window[11][7];
assign temp[1128] = ~window[11][8];
assign temp[1152] = window[12][0];
assign temp[1153] = window[12][1];
assign temp[1154] = window[12][2];
assign temp[1155] = ~window[12][3];
assign temp[1156] = ~window[12][4];
assign temp[1157] = ~window[12][5];
assign temp[1158] = ~window[12][6];
assign temp[1159] = window[12][7];
assign temp[1160] = window[12][8];
assign temp[1184] = window[13][0];
assign temp[1185] = window[13][1];
assign temp[1186] = window[13][2];
assign temp[1187] = window[13][3];
assign temp[1188] = window[13][4];
assign temp[1189] = window[13][5];
assign temp[1190] = ~window[13][6];
assign temp[1191] = ~window[13][7];
assign temp[1192] = window[13][8];
assign temp[1216] = ~window[14][0];
assign temp[1217] = ~window[14][1];
assign temp[1218] = ~window[14][2];
assign temp[1219] = window[14][3];
assign temp[1220] = ~window[14][4];
assign temp[1221] = ~window[14][5];
assign temp[1222] = window[14][6];
assign temp[1223] = ~window[14][7];
assign temp[1224] = ~window[14][8];
assign temp[1248] = window[15][0];
assign temp[1249] = window[15][1];
assign temp[1250] = window[15][2];
assign temp[1251] = ~window[15][3];
assign temp[1252] = window[15][4];
assign temp[1253] = ~window[15][5];
assign temp[1254] = window[15][6];
assign temp[1255] = window[15][7];
assign temp[1256] = ~window[15][8];
assign temp[1280] = ~window[16][0];
assign temp[1281] = window[16][1];
assign temp[1282] = window[16][2];
assign temp[1283] = ~window[16][3];
assign temp[1284] = window[16][4];
assign temp[1285] = window[16][5];
assign temp[1286] = ~window[16][6];
assign temp[1287] = ~window[16][7];
assign temp[1288] = window[16][8];
assign temp[1312] = window[17][0];
assign temp[1313] = ~window[17][1];
assign temp[1314] = ~window[17][2];
assign temp[1315] = window[17][3];
assign temp[1316] = window[17][4];
assign temp[1317] = window[17][5];
assign temp[1318] = window[17][6];
assign temp[1319] = window[17][7];
assign temp[1320] = window[17][8];
assign temp[1344] = ~window[18][0];
assign temp[1345] = ~window[18][1];
assign temp[1346] = ~window[18][2];
assign temp[1347] = ~window[18][3];
assign temp[1348] = window[18][4];
assign temp[1349] = window[18][5];
assign temp[1350] = window[18][6];
assign temp[1351] = window[18][7];
assign temp[1352] = ~window[18][8];
assign temp[1376] = window[19][0];
assign temp[1377] = ~window[19][1];
assign temp[1378] = window[19][2];
assign temp[1379] = window[19][3];
assign temp[1380] = ~window[19][4];
assign temp[1381] = ~window[19][5];
assign temp[1382] = window[19][6];
assign temp[1383] = window[19][7];
assign temp[1384] = ~window[19][8];
assign temp[1408] = window[20][0];
assign temp[1409] = ~window[20][1];
assign temp[1410] = ~window[20][2];
assign temp[1411] = ~window[20][3];
assign temp[1412] = window[20][4];
assign temp[1413] = window[20][5];
assign temp[1414] = window[20][6];
assign temp[1415] = ~window[20][7];
assign temp[1416] = window[20][8];
assign temp[1440] = window[21][0];
assign temp[1441] = ~window[21][1];
assign temp[1442] = ~window[21][2];
assign temp[1443] = window[21][3];
assign temp[1444] = ~window[21][4];
assign temp[1445] = window[21][5];
assign temp[1446] = window[21][6];
assign temp[1447] = window[21][7];
assign temp[1448] = ~window[21][8];
assign temp[1472] = window[22][0];
assign temp[1473] = window[22][1];
assign temp[1474] = window[22][2];
assign temp[1475] = window[22][3];
assign temp[1476] = ~window[22][4];
assign temp[1477] = ~window[22][5];
assign temp[1478] = window[22][6];
assign temp[1479] = ~window[22][7];
assign temp[1480] = window[22][8];
assign temp[1504] = ~window[23][0];
assign temp[1505] = ~window[23][1];
assign temp[1506] = ~window[23][2];
assign temp[1507] = window[23][3];
assign temp[1508] = ~window[23][4];
assign temp[1509] = ~window[23][5];
assign temp[1510] = ~window[23][6];
assign temp[1511] = ~window[23][7];
assign temp[1512] = ~window[23][8];
assign temp[1536] = ~window[24][0];
assign temp[1537] = ~window[24][1];
assign temp[1538] = ~window[24][2];
assign temp[1539] = window[24][3];
assign temp[1540] = ~window[24][4];
assign temp[1541] = ~window[24][5];
assign temp[1542] = ~window[24][6];
assign temp[1543] = window[24][7];
assign temp[1544] = window[24][8];
assign temp[1568] = window[25][0];
assign temp[1569] = ~window[25][1];
assign temp[1570] = ~window[25][2];
assign temp[1571] = window[25][3];
assign temp[1572] = window[25][4];
assign temp[1573] = window[25][5];
assign temp[1574] = window[25][6];
assign temp[1575] = ~window[25][7];
assign temp[1576] = window[25][8];
assign temp[1600] = window[26][0];
assign temp[1601] = ~window[26][1];
assign temp[1602] = ~window[26][2];
assign temp[1603] = window[26][3];
assign temp[1604] = window[26][4];
assign temp[1605] = ~window[26][5];
assign temp[1606] = window[26][6];
assign temp[1607] = window[26][7];
assign temp[1608] = window[26][8];
assign temp[1632] = window[27][0];
assign temp[1633] = window[27][1];
assign temp[1634] = window[27][2];
assign temp[1635] = window[27][3];
assign temp[1636] = window[27][4];
assign temp[1637] = window[27][5];
assign temp[1638] = window[27][6];
assign temp[1639] = ~window[27][7];
assign temp[1640] = ~window[27][8];
assign temp[1664] = ~window[28][0];
assign temp[1665] = window[28][1];
assign temp[1666] = window[28][2];
assign temp[1667] = ~window[28][3];
assign temp[1668] = window[28][4];
assign temp[1669] = window[28][5];
assign temp[1670] = ~window[28][6];
assign temp[1671] = ~window[28][7];
assign temp[1672] = window[28][8];
assign temp[1696] = window[29][0];
assign temp[1697] = window[29][1];
assign temp[1698] = window[29][2];
assign temp[1699] = window[29][3];
assign temp[1700] = window[29][4];
assign temp[1701] = window[29][5];
assign temp[1702] = window[29][6];
assign temp[1703] = ~window[29][7];
assign temp[1704] = window[29][8];
assign temp[1728] = ~window[30][0];
assign temp[1729] = ~window[30][1];
assign temp[1730] = window[30][2];
assign temp[1731] = ~window[30][3];
assign temp[1732] = ~window[30][4];
assign temp[1733] = window[30][5];
assign temp[1734] = ~window[30][6];
assign temp[1735] = ~window[30][7];
assign temp[1736] = window[30][8];
assign temp[1760] = ~window[31][0];
assign temp[1761] = ~window[31][1];
assign temp[1762] = ~window[31][2];
assign temp[1763] = ~window[31][3];
assign temp[1764] = ~window[31][4];
assign temp[1765] = window[31][5];
assign temp[1766] = ~window[31][6];
assign temp[1767] = window[31][7];
assign temp[1768] = window[31][8];
assign temp[800] = ~window[0][0];
assign temp[801] = window[0][1];
assign temp[802] = window[0][2];
assign temp[803] = window[0][3];
assign temp[804] = window[0][4];
assign temp[805] = window[0][5];
assign temp[806] = window[0][6];
assign temp[807] = window[0][7];
assign temp[808] = window[0][8];
assign temp[832] = ~window[1][0];
assign temp[833] = window[1][1];
assign temp[834] = window[1][2];
assign temp[835] = ~window[1][3];
assign temp[836] = ~window[1][4];
assign temp[837] = ~window[1][5];
assign temp[838] = window[1][6];
assign temp[839] = window[1][7];
assign temp[840] = ~window[1][8];
assign temp[864] = window[2][0];
assign temp[865] = window[2][1];
assign temp[866] = window[2][2];
assign temp[867] = window[2][3];
assign temp[868] = ~window[2][4];
assign temp[869] = ~window[2][5];
assign temp[870] = window[2][6];
assign temp[871] = window[2][7];
assign temp[872] = window[2][8];
assign temp[896] = window[3][0];
assign temp[897] = ~window[3][1];
assign temp[898] = window[3][2];
assign temp[899] = window[3][3];
assign temp[900] = window[3][4];
assign temp[901] = ~window[3][5];
assign temp[902] = window[3][6];
assign temp[903] = window[3][7];
assign temp[904] = window[3][8];
assign temp[928] = window[4][0];
assign temp[929] = window[4][1];
assign temp[930] = ~window[4][2];
assign temp[931] = window[4][3];
assign temp[932] = window[4][4];
assign temp[933] = window[4][5];
assign temp[934] = window[4][6];
assign temp[935] = window[4][7];
assign temp[936] = window[4][8];
assign temp[960] = ~window[5][0];
assign temp[961] = ~window[5][1];
assign temp[962] = ~window[5][2];
assign temp[963] = window[5][3];
assign temp[964] = ~window[5][4];
assign temp[965] = window[5][5];
assign temp[966] = window[5][6];
assign temp[967] = ~window[5][7];
assign temp[968] = window[5][8];
assign temp[992] = ~window[6][0];
assign temp[993] = ~window[6][1];
assign temp[994] = ~window[6][2];
assign temp[995] = window[6][3];
assign temp[996] = window[6][4];
assign temp[997] = window[6][5];
assign temp[998] = window[6][6];
assign temp[999] = window[6][7];
assign temp[1000] = window[6][8];
assign temp[1024] = ~window[7][0];
assign temp[1025] = window[7][1];
assign temp[1026] = ~window[7][2];
assign temp[1027] = ~window[7][3];
assign temp[1028] = ~window[7][4];
assign temp[1029] = window[7][5];
assign temp[1030] = window[7][6];
assign temp[1031] = window[7][7];
assign temp[1032] = window[7][8];
assign temp[1056] = ~window[8][0];
assign temp[1057] = window[8][1];
assign temp[1058] = ~window[8][2];
assign temp[1059] = window[8][3];
assign temp[1060] = window[8][4];
assign temp[1061] = window[8][5];
assign temp[1062] = window[8][6];
assign temp[1063] = window[8][7];
assign temp[1064] = window[8][8];
assign temp[1088] = window[9][0];
assign temp[1089] = window[9][1];
assign temp[1090] = ~window[9][2];
assign temp[1091] = window[9][3];
assign temp[1092] = ~window[9][4];
assign temp[1093] = ~window[9][5];
assign temp[1094] = window[9][6];
assign temp[1095] = window[9][7];
assign temp[1096] = window[9][8];
assign temp[1120] = window[10][0];
assign temp[1121] = window[10][1];
assign temp[1122] = window[10][2];
assign temp[1123] = window[10][3];
assign temp[1124] = ~window[10][4];
assign temp[1125] = window[10][5];
assign temp[1126] = window[10][6];
assign temp[1127] = ~window[10][7];
assign temp[1128] = ~window[10][8];
assign temp[1152] = window[11][0];
assign temp[1153] = window[11][1];
assign temp[1154] = window[11][2];
assign temp[1155] = window[11][3];
assign temp[1156] = ~window[11][4];
assign temp[1157] = window[11][5];
assign temp[1158] = window[11][6];
assign temp[1159] = ~window[11][7];
assign temp[1160] = ~window[11][8];
assign temp[1184] = window[12][0];
assign temp[1185] = window[12][1];
assign temp[1186] = window[12][2];
assign temp[1187] = window[12][3];
assign temp[1188] = ~window[12][4];
assign temp[1189] = ~window[12][5];
assign temp[1190] = ~window[12][6];
assign temp[1191] = ~window[12][7];
assign temp[1192] = window[12][8];
assign temp[1216] = window[13][0];
assign temp[1217] = ~window[13][1];
assign temp[1218] = window[13][2];
assign temp[1219] = window[13][3];
assign temp[1220] = ~window[13][4];
assign temp[1221] = window[13][5];
assign temp[1222] = ~window[13][6];
assign temp[1223] = ~window[13][7];
assign temp[1224] = ~window[13][8];
assign temp[1248] = ~window[14][0];
assign temp[1249] = window[14][1];
assign temp[1250] = ~window[14][2];
assign temp[1251] = window[14][3];
assign temp[1252] = ~window[14][4];
assign temp[1253] = window[14][5];
assign temp[1254] = window[14][6];
assign temp[1255] = ~window[14][7];
assign temp[1256] = window[14][8];
assign temp[1280] = window[15][0];
assign temp[1281] = window[15][1];
assign temp[1282] = window[15][2];
assign temp[1283] = ~window[15][3];
assign temp[1284] = window[15][4];
assign temp[1285] = ~window[15][5];
assign temp[1286] = window[15][6];
assign temp[1287] = window[15][7];
assign temp[1288] = ~window[15][8];
assign temp[1312] = window[16][0];
assign temp[1313] = ~window[16][1];
assign temp[1314] = ~window[16][2];
assign temp[1315] = ~window[16][3];
assign temp[1316] = window[16][4];
assign temp[1317] = window[16][5];
assign temp[1318] = ~window[16][6];
assign temp[1319] = window[16][7];
assign temp[1320] = ~window[16][8];
assign temp[1344] = window[17][0];
assign temp[1345] = window[17][1];
assign temp[1346] = window[17][2];
assign temp[1347] = ~window[17][3];
assign temp[1348] = ~window[17][4];
assign temp[1349] = ~window[17][5];
assign temp[1350] = window[17][6];
assign temp[1351] = window[17][7];
assign temp[1352] = window[17][8];
assign temp[1376] = ~window[18][0];
assign temp[1377] = window[18][1];
assign temp[1378] = window[18][2];
assign temp[1379] = window[18][3];
assign temp[1380] = ~window[18][4];
assign temp[1381] = window[18][5];
assign temp[1382] = window[18][6];
assign temp[1383] = window[18][7];
assign temp[1384] = window[18][8];
assign temp[1408] = ~window[19][0];
assign temp[1409] = ~window[19][1];
assign temp[1410] = window[19][2];
assign temp[1411] = ~window[19][3];
assign temp[1412] = ~window[19][4];
assign temp[1413] = ~window[19][5];
assign temp[1414] = ~window[19][6];
assign temp[1415] = ~window[19][7];
assign temp[1416] = ~window[19][8];
assign temp[1440] = window[20][0];
assign temp[1441] = window[20][1];
assign temp[1442] = window[20][2];
assign temp[1443] = window[20][3];
assign temp[1444] = window[20][4];
assign temp[1445] = ~window[20][5];
assign temp[1446] = ~window[20][6];
assign temp[1447] = window[20][7];
assign temp[1448] = window[20][8];
assign temp[1472] = ~window[21][0];
assign temp[1473] = window[21][1];
assign temp[1474] = ~window[21][2];
assign temp[1475] = ~window[21][3];
assign temp[1476] = ~window[21][4];
assign temp[1477] = ~window[21][5];
assign temp[1478] = window[21][6];
assign temp[1479] = ~window[21][7];
assign temp[1480] = ~window[21][8];
assign temp[1504] = window[22][0];
assign temp[1505] = ~window[22][1];
assign temp[1506] = window[22][2];
assign temp[1507] = ~window[22][3];
assign temp[1508] = window[22][4];
assign temp[1509] = window[22][5];
assign temp[1510] = window[22][6];
assign temp[1511] = ~window[22][7];
assign temp[1512] = ~window[22][8];
assign temp[1536] = ~window[23][0];
assign temp[1537] = window[23][1];
assign temp[1538] = ~window[23][2];
assign temp[1539] = window[23][3];
assign temp[1540] = ~window[23][4];
assign temp[1541] = ~window[23][5];
assign temp[1542] = window[23][6];
assign temp[1543] = window[23][7];
assign temp[1544] = window[23][8];
assign temp[1568] = window[24][0];
assign temp[1569] = window[24][1];
assign temp[1570] = window[24][2];
assign temp[1571] = window[24][3];
assign temp[1572] = ~window[24][4];
assign temp[1573] = ~window[24][5];
assign temp[1574] = window[24][6];
assign temp[1575] = window[24][7];
assign temp[1576] = window[24][8];
assign temp[1600] = window[25][0];
assign temp[1601] = window[25][1];
assign temp[1602] = ~window[25][2];
assign temp[1603] = ~window[25][3];
assign temp[1604] = window[25][4];
assign temp[1605] = window[25][5];
assign temp[1606] = ~window[25][6];
assign temp[1607] = window[25][7];
assign temp[1608] = window[25][8];
assign temp[1632] = ~window[26][0];
assign temp[1633] = window[26][1];
assign temp[1634] = window[26][2];
assign temp[1635] = ~window[26][3];
assign temp[1636] = ~window[26][4];
assign temp[1637] = ~window[26][5];
assign temp[1638] = ~window[26][6];
assign temp[1639] = ~window[26][7];
assign temp[1640] = ~window[26][8];
assign temp[1664] = ~window[27][0];
assign temp[1665] = ~window[27][1];
assign temp[1666] = ~window[27][2];
assign temp[1667] = ~window[27][3];
assign temp[1668] = window[27][4];
assign temp[1669] = window[27][5];
assign temp[1670] = window[27][6];
assign temp[1671] = ~window[27][7];
assign temp[1672] = window[27][8];
assign temp[1696] = window[28][0];
assign temp[1697] = ~window[28][1];
assign temp[1698] = window[28][2];
assign temp[1699] = window[28][3];
assign temp[1700] = window[28][4];
assign temp[1701] = window[28][5];
assign temp[1702] = ~window[28][6];
assign temp[1703] = ~window[28][7];
assign temp[1704] = ~window[28][8];
assign temp[1728] = window[29][0];
assign temp[1729] = window[29][1];
assign temp[1730] = window[29][2];
assign temp[1731] = ~window[29][3];
assign temp[1732] = window[29][4];
assign temp[1733] = window[29][5];
assign temp[1734] = window[29][6];
assign temp[1735] = ~window[29][7];
assign temp[1736] = ~window[29][8];
assign temp[1760] = ~window[30][0];
assign temp[1761] = ~window[30][1];
assign temp[1762] = ~window[30][2];
assign temp[1763] = ~window[30][3];
assign temp[1764] = ~window[30][4];
assign temp[1765] = window[30][5];
assign temp[1766] = ~window[30][6];
assign temp[1767] = ~window[30][7];
assign temp[1768] = ~window[30][8];
assign temp[1792] = window[31][0];
assign temp[1793] = window[31][1];
assign temp[1794] = window[31][2];
assign temp[1795] = window[31][3];
assign temp[1796] = ~window[31][4];
assign temp[1797] = ~window[31][5];
assign temp[1798] = ~window[31][6];
assign temp[1799] = window[31][7];
assign temp[1800] = window[31][8];
assign temp[832] = ~window[0][0];
assign temp[833] = ~window[0][1];
assign temp[834] = window[0][2];
assign temp[835] = ~window[0][3];
assign temp[836] = ~window[0][4];
assign temp[837] = window[0][5];
assign temp[838] = window[0][6];
assign temp[839] = ~window[0][7];
assign temp[840] = window[0][8];
assign temp[864] = window[1][0];
assign temp[865] = ~window[1][1];
assign temp[866] = ~window[1][2];
assign temp[867] = window[1][3];
assign temp[868] = window[1][4];
assign temp[869] = window[1][5];
assign temp[870] = window[1][6];
assign temp[871] = ~window[1][7];
assign temp[872] = window[1][8];
assign temp[896] = ~window[2][0];
assign temp[897] = ~window[2][1];
assign temp[898] = ~window[2][2];
assign temp[899] = window[2][3];
assign temp[900] = ~window[2][4];
assign temp[901] = window[2][5];
assign temp[902] = ~window[2][6];
assign temp[903] = window[2][7];
assign temp[904] = window[2][8];
assign temp[928] = ~window[3][0];
assign temp[929] = ~window[3][1];
assign temp[930] = ~window[3][2];
assign temp[931] = ~window[3][3];
assign temp[932] = ~window[3][4];
assign temp[933] = window[3][5];
assign temp[934] = ~window[3][6];
assign temp[935] = ~window[3][7];
assign temp[936] = window[3][8];
assign temp[960] = ~window[4][0];
assign temp[961] = ~window[4][1];
assign temp[962] = ~window[4][2];
assign temp[963] = ~window[4][3];
assign temp[964] = ~window[4][4];
assign temp[965] = ~window[4][5];
assign temp[966] = ~window[4][6];
assign temp[967] = ~window[4][7];
assign temp[968] = window[4][8];
assign temp[992] = ~window[5][0];
assign temp[993] = window[5][1];
assign temp[994] = window[5][2];
assign temp[995] = window[5][3];
assign temp[996] = window[5][4];
assign temp[997] = window[5][5];
assign temp[998] = ~window[5][6];
assign temp[999] = window[5][7];
assign temp[1000] = window[5][8];
assign temp[1024] = ~window[6][0];
assign temp[1025] = window[6][1];
assign temp[1026] = ~window[6][2];
assign temp[1027] = ~window[6][3];
assign temp[1028] = ~window[6][4];
assign temp[1029] = ~window[6][5];
assign temp[1030] = window[6][6];
assign temp[1031] = window[6][7];
assign temp[1032] = ~window[6][8];
assign temp[1056] = ~window[7][0];
assign temp[1057] = ~window[7][1];
assign temp[1058] = window[7][2];
assign temp[1059] = ~window[7][3];
assign temp[1060] = ~window[7][4];
assign temp[1061] = window[7][5];
assign temp[1062] = ~window[7][6];
assign temp[1063] = ~window[7][7];
assign temp[1064] = window[7][8];
assign temp[1088] = ~window[8][0];
assign temp[1089] = ~window[8][1];
assign temp[1090] = window[8][2];
assign temp[1091] = ~window[8][3];
assign temp[1092] = ~window[8][4];
assign temp[1093] = window[8][5];
assign temp[1094] = ~window[8][6];
assign temp[1095] = ~window[8][7];
assign temp[1096] = ~window[8][8];
assign temp[1120] = ~window[9][0];
assign temp[1121] = ~window[9][1];
assign temp[1122] = window[9][2];
assign temp[1123] = ~window[9][3];
assign temp[1124] = ~window[9][4];
assign temp[1125] = window[9][5];
assign temp[1126] = ~window[9][6];
assign temp[1127] = ~window[9][7];
assign temp[1128] = window[9][8];
assign temp[1152] = ~window[10][0];
assign temp[1153] = ~window[10][1];
assign temp[1154] = ~window[10][2];
assign temp[1155] = ~window[10][3];
assign temp[1156] = ~window[10][4];
assign temp[1157] = window[10][5];
assign temp[1158] = ~window[10][6];
assign temp[1159] = ~window[10][7];
assign temp[1160] = ~window[10][8];
assign temp[1184] = window[11][0];
assign temp[1185] = window[11][1];
assign temp[1186] = ~window[11][2];
assign temp[1187] = window[11][3];
assign temp[1188] = ~window[11][4];
assign temp[1189] = window[11][5];
assign temp[1190] = window[11][6];
assign temp[1191] = ~window[11][7];
assign temp[1192] = ~window[11][8];
assign temp[1216] = window[12][0];
assign temp[1217] = window[12][1];
assign temp[1218] = ~window[12][2];
assign temp[1219] = ~window[12][3];
assign temp[1220] = ~window[12][4];
assign temp[1221] = ~window[12][5];
assign temp[1222] = window[12][6];
assign temp[1223] = window[12][7];
assign temp[1224] = window[12][8];
assign temp[1248] = window[13][0];
assign temp[1249] = window[13][1];
assign temp[1250] = ~window[13][2];
assign temp[1251] = window[13][3];
assign temp[1252] = window[13][4];
assign temp[1253] = window[13][5];
assign temp[1254] = window[13][6];
assign temp[1255] = ~window[13][7];
assign temp[1256] = ~window[13][8];
assign temp[1280] = window[14][0];
assign temp[1281] = ~window[14][1];
assign temp[1282] = ~window[14][2];
assign temp[1283] = ~window[14][3];
assign temp[1284] = ~window[14][4];
assign temp[1285] = ~window[14][5];
assign temp[1286] = ~window[14][6];
assign temp[1287] = ~window[14][7];
assign temp[1288] = ~window[14][8];
assign temp[1312] = ~window[15][0];
assign temp[1313] = window[15][1];
assign temp[1314] = ~window[15][2];
assign temp[1315] = ~window[15][3];
assign temp[1316] = window[15][4];
assign temp[1317] = ~window[15][5];
assign temp[1318] = ~window[15][6];
assign temp[1319] = window[15][7];
assign temp[1320] = ~window[15][8];
assign temp[1344] = ~window[16][0];
assign temp[1345] = window[16][1];
assign temp[1346] = window[16][2];
assign temp[1347] = ~window[16][3];
assign temp[1348] = window[16][4];
assign temp[1349] = window[16][5];
assign temp[1350] = ~window[16][6];
assign temp[1351] = ~window[16][7];
assign temp[1352] = ~window[16][8];
assign temp[1376] = window[17][0];
assign temp[1377] = ~window[17][1];
assign temp[1378] = window[17][2];
assign temp[1379] = ~window[17][3];
assign temp[1380] = ~window[17][4];
assign temp[1381] = window[17][5];
assign temp[1382] = ~window[17][6];
assign temp[1383] = ~window[17][7];
assign temp[1384] = window[17][8];
assign temp[1408] = ~window[18][0];
assign temp[1409] = window[18][1];
assign temp[1410] = ~window[18][2];
assign temp[1411] = window[18][3];
assign temp[1412] = window[18][4];
assign temp[1413] = ~window[18][5];
assign temp[1414] = ~window[18][6];
assign temp[1415] = window[18][7];
assign temp[1416] = window[18][8];
assign temp[1440] = window[19][0];
assign temp[1441] = window[19][1];
assign temp[1442] = ~window[19][2];
assign temp[1443] = window[19][3];
assign temp[1444] = ~window[19][4];
assign temp[1445] = window[19][5];
assign temp[1446] = window[19][6];
assign temp[1447] = ~window[19][7];
assign temp[1448] = window[19][8];
assign temp[1472] = ~window[20][0];
assign temp[1473] = ~window[20][1];
assign temp[1474] = ~window[20][2];
assign temp[1475] = ~window[20][3];
assign temp[1476] = ~window[20][4];
assign temp[1477] = window[20][5];
assign temp[1478] = ~window[20][6];
assign temp[1479] = ~window[20][7];
assign temp[1480] = window[20][8];
assign temp[1504] = ~window[21][0];
assign temp[1505] = window[21][1];
assign temp[1506] = ~window[21][2];
assign temp[1507] = window[21][3];
assign temp[1508] = window[21][4];
assign temp[1509] = window[21][5];
assign temp[1510] = window[21][6];
assign temp[1511] = window[21][7];
assign temp[1512] = window[21][8];
assign temp[1536] = window[22][0];
assign temp[1537] = window[22][1];
assign temp[1538] = window[22][2];
assign temp[1539] = window[22][3];
assign temp[1540] = window[22][4];
assign temp[1541] = ~window[22][5];
assign temp[1542] = window[22][6];
assign temp[1543] = ~window[22][7];
assign temp[1544] = ~window[22][8];
assign temp[1568] = ~window[23][0];
assign temp[1569] = window[23][1];
assign temp[1570] = ~window[23][2];
assign temp[1571] = ~window[23][3];
assign temp[1572] = ~window[23][4];
assign temp[1573] = window[23][5];
assign temp[1574] = window[23][6];
assign temp[1575] = ~window[23][7];
assign temp[1576] = window[23][8];
assign temp[1600] = window[24][0];
assign temp[1601] = ~window[24][1];
assign temp[1602] = ~window[24][2];
assign temp[1603] = window[24][3];
assign temp[1604] = ~window[24][4];
assign temp[1605] = ~window[24][5];
assign temp[1606] = ~window[24][6];
assign temp[1607] = window[24][7];
assign temp[1608] = window[24][8];
assign temp[1632] = ~window[25][0];
assign temp[1633] = window[25][1];
assign temp[1634] = window[25][2];
assign temp[1635] = ~window[25][3];
assign temp[1636] = window[25][4];
assign temp[1637] = ~window[25][5];
assign temp[1638] = ~window[25][6];
assign temp[1639] = window[25][7];
assign temp[1640] = ~window[25][8];
assign temp[1664] = window[26][0];
assign temp[1665] = window[26][1];
assign temp[1666] = ~window[26][2];
assign temp[1667] = window[26][3];
assign temp[1668] = ~window[26][4];
assign temp[1669] = window[26][5];
assign temp[1670] = window[26][6];
assign temp[1671] = ~window[26][7];
assign temp[1672] = window[26][8];
assign temp[1696] = ~window[27][0];
assign temp[1697] = ~window[27][1];
assign temp[1698] = window[27][2];
assign temp[1699] = ~window[27][3];
assign temp[1700] = ~window[27][4];
assign temp[1701] = window[27][5];
assign temp[1702] = ~window[27][6];
assign temp[1703] = ~window[27][7];
assign temp[1704] = ~window[27][8];
assign temp[1728] = ~window[28][0];
assign temp[1729] = window[28][1];
assign temp[1730] = ~window[28][2];
assign temp[1731] = window[28][3];
assign temp[1732] = window[28][4];
assign temp[1733] = ~window[28][5];
assign temp[1734] = ~window[28][6];
assign temp[1735] = ~window[28][7];
assign temp[1736] = ~window[28][8];
assign temp[1760] = window[29][0];
assign temp[1761] = window[29][1];
assign temp[1762] = window[29][2];
assign temp[1763] = window[29][3];
assign temp[1764] = ~window[29][4];
assign temp[1765] = window[29][5];
assign temp[1766] = ~window[29][6];
assign temp[1767] = ~window[29][7];
assign temp[1768] = ~window[29][8];
assign temp[1792] = window[30][0];
assign temp[1793] = window[30][1];
assign temp[1794] = window[30][2];
assign temp[1795] = window[30][3];
assign temp[1796] = window[30][4];
assign temp[1797] = window[30][5];
assign temp[1798] = window[30][6];
assign temp[1799] = window[30][7];
assign temp[1800] = window[30][8];
assign temp[1824] = window[31][0];
assign temp[1825] = window[31][1];
assign temp[1826] = ~window[31][2];
assign temp[1827] = window[31][3];
assign temp[1828] = ~window[31][4];
assign temp[1829] = window[31][5];
assign temp[1830] = ~window[31][6];
assign temp[1831] = ~window[31][7];
assign temp[1832] = ~window[31][8];
assign temp[864] = ~window[0][0];
assign temp[865] = window[0][1];
assign temp[866] = ~window[0][2];
assign temp[867] = window[0][3];
assign temp[868] = window[0][4];
assign temp[869] = window[0][5];
assign temp[870] = window[0][6];
assign temp[871] = window[0][7];
assign temp[872] = window[0][8];
assign temp[896] = ~window[1][0];
assign temp[897] = window[1][1];
assign temp[898] = window[1][2];
assign temp[899] = window[1][3];
assign temp[900] = ~window[1][4];
assign temp[901] = window[1][5];
assign temp[902] = window[1][6];
assign temp[903] = ~window[1][7];
assign temp[904] = ~window[1][8];
assign temp[928] = ~window[2][0];
assign temp[929] = ~window[2][1];
assign temp[930] = ~window[2][2];
assign temp[931] = window[2][3];
assign temp[932] = ~window[2][4];
assign temp[933] = ~window[2][5];
assign temp[934] = ~window[2][6];
assign temp[935] = window[2][7];
assign temp[936] = ~window[2][8];
assign temp[960] = window[3][0];
assign temp[961] = ~window[3][1];
assign temp[962] = ~window[3][2];
assign temp[963] = window[3][3];
assign temp[964] = ~window[3][4];
assign temp[965] = ~window[3][5];
assign temp[966] = window[3][6];
assign temp[967] = window[3][7];
assign temp[968] = ~window[3][8];
assign temp[992] = window[4][0];
assign temp[993] = window[4][1];
assign temp[994] = window[4][2];
assign temp[995] = ~window[4][3];
assign temp[996] = window[4][4];
assign temp[997] = window[4][5];
assign temp[998] = window[4][6];
assign temp[999] = ~window[4][7];
assign temp[1000] = window[4][8];
assign temp[1024] = window[5][0];
assign temp[1025] = ~window[5][1];
assign temp[1026] = ~window[5][2];
assign temp[1027] = window[5][3];
assign temp[1028] = window[5][4];
assign temp[1029] = window[5][5];
assign temp[1030] = window[5][6];
assign temp[1031] = window[5][7];
assign temp[1032] = window[5][8];
assign temp[1056] = ~window[6][0];
assign temp[1057] = window[6][1];
assign temp[1058] = ~window[6][2];
assign temp[1059] = ~window[6][3];
assign temp[1060] = ~window[6][4];
assign temp[1061] = window[6][5];
assign temp[1062] = window[6][6];
assign temp[1063] = window[6][7];
assign temp[1064] = window[6][8];
assign temp[1088] = window[7][0];
assign temp[1089] = window[7][1];
assign temp[1090] = ~window[7][2];
assign temp[1091] = window[7][3];
assign temp[1092] = window[7][4];
assign temp[1093] = window[7][5];
assign temp[1094] = ~window[7][6];
assign temp[1095] = window[7][7];
assign temp[1096] = window[7][8];
assign temp[1120] = ~window[8][0];
assign temp[1121] = window[8][1];
assign temp[1122] = ~window[8][2];
assign temp[1123] = window[8][3];
assign temp[1124] = window[8][4];
assign temp[1125] = ~window[8][5];
assign temp[1126] = window[8][6];
assign temp[1127] = window[8][7];
assign temp[1128] = window[8][8];
assign temp[1152] = window[9][0];
assign temp[1153] = window[9][1];
assign temp[1154] = ~window[9][2];
assign temp[1155] = ~window[9][3];
assign temp[1156] = window[9][4];
assign temp[1157] = ~window[9][5];
assign temp[1158] = window[9][6];
assign temp[1159] = window[9][7];
assign temp[1160] = window[9][8];
assign temp[1184] = window[10][0];
assign temp[1185] = window[10][1];
assign temp[1186] = ~window[10][2];
assign temp[1187] = window[10][3];
assign temp[1188] = window[10][4];
assign temp[1189] = window[10][5];
assign temp[1190] = window[10][6];
assign temp[1191] = ~window[10][7];
assign temp[1192] = window[10][8];
assign temp[1216] = ~window[11][0];
assign temp[1217] = window[11][1];
assign temp[1218] = window[11][2];
assign temp[1219] = ~window[11][3];
assign temp[1220] = window[11][4];
assign temp[1221] = window[11][5];
assign temp[1222] = ~window[11][6];
assign temp[1223] = ~window[11][7];
assign temp[1224] = window[11][8];
assign temp[1248] = ~window[12][0];
assign temp[1249] = window[12][1];
assign temp[1250] = window[12][2];
assign temp[1251] = ~window[12][3];
assign temp[1252] = ~window[12][4];
assign temp[1253] = ~window[12][5];
assign temp[1254] = ~window[12][6];
assign temp[1255] = ~window[12][7];
assign temp[1256] = ~window[12][8];
assign temp[1280] = ~window[13][0];
assign temp[1281] = window[13][1];
assign temp[1282] = ~window[13][2];
assign temp[1283] = ~window[13][3];
assign temp[1284] = ~window[13][4];
assign temp[1285] = ~window[13][5];
assign temp[1286] = ~window[13][6];
assign temp[1287] = ~window[13][7];
assign temp[1288] = ~window[13][8];
assign temp[1312] = window[14][0];
assign temp[1313] = ~window[14][1];
assign temp[1314] = ~window[14][2];
assign temp[1315] = window[14][3];
assign temp[1316] = ~window[14][4];
assign temp[1317] = ~window[14][5];
assign temp[1318] = window[14][6];
assign temp[1319] = window[14][7];
assign temp[1320] = ~window[14][8];
assign temp[1344] = window[15][0];
assign temp[1345] = ~window[15][1];
assign temp[1346] = window[15][2];
assign temp[1347] = window[15][3];
assign temp[1348] = window[15][4];
assign temp[1349] = window[15][5];
assign temp[1350] = window[15][6];
assign temp[1351] = window[15][7];
assign temp[1352] = window[15][8];
assign temp[1376] = window[16][0];
assign temp[1377] = ~window[16][1];
assign temp[1378] = ~window[16][2];
assign temp[1379] = ~window[16][3];
assign temp[1380] = window[16][4];
assign temp[1381] = window[16][5];
assign temp[1382] = ~window[16][6];
assign temp[1383] = window[16][7];
assign temp[1384] = window[16][8];
assign temp[1408] = window[17][0];
assign temp[1409] = window[17][1];
assign temp[1410] = window[17][2];
assign temp[1411] = window[17][3];
assign temp[1412] = ~window[17][4];
assign temp[1413] = ~window[17][5];
assign temp[1414] = ~window[17][6];
assign temp[1415] = ~window[17][7];
assign temp[1416] = window[17][8];
assign temp[1440] = window[18][0];
assign temp[1441] = ~window[18][1];
assign temp[1442] = ~window[18][2];
assign temp[1443] = window[18][3];
assign temp[1444] = window[18][4];
assign temp[1445] = ~window[18][5];
assign temp[1446] = ~window[18][6];
assign temp[1447] = window[18][7];
assign temp[1448] = ~window[18][8];
assign temp[1472] = window[19][0];
assign temp[1473] = ~window[19][1];
assign temp[1474] = window[19][2];
assign temp[1475] = ~window[19][3];
assign temp[1476] = ~window[19][4];
assign temp[1477] = window[19][5];
assign temp[1478] = window[19][6];
assign temp[1479] = ~window[19][7];
assign temp[1480] = ~window[19][8];
assign temp[1504] = ~window[20][0];
assign temp[1505] = ~window[20][1];
assign temp[1506] = ~window[20][2];
assign temp[1507] = window[20][3];
assign temp[1508] = ~window[20][4];
assign temp[1509] = ~window[20][5];
assign temp[1510] = window[20][6];
assign temp[1511] = ~window[20][7];
assign temp[1512] = window[20][8];
assign temp[1536] = window[21][0];
assign temp[1537] = window[21][1];
assign temp[1538] = window[21][2];
assign temp[1539] = window[21][3];
assign temp[1540] = window[21][4];
assign temp[1541] = window[21][5];
assign temp[1542] = window[21][6];
assign temp[1543] = ~window[21][7];
assign temp[1544] = window[21][8];
assign temp[1568] = ~window[22][0];
assign temp[1569] = window[22][1];
assign temp[1570] = window[22][2];
assign temp[1571] = ~window[22][3];
assign temp[1572] = ~window[22][4];
assign temp[1573] = window[22][5];
assign temp[1574] = ~window[22][6];
assign temp[1575] = ~window[22][7];
assign temp[1576] = ~window[22][8];
assign temp[1600] = window[23][0];
assign temp[1601] = ~window[23][1];
assign temp[1602] = ~window[23][2];
assign temp[1603] = window[23][3];
assign temp[1604] = window[23][4];
assign temp[1605] = ~window[23][5];
assign temp[1606] = window[23][6];
assign temp[1607] = window[23][7];
assign temp[1608] = ~window[23][8];
assign temp[1632] = ~window[24][0];
assign temp[1633] = ~window[24][1];
assign temp[1634] = ~window[24][2];
assign temp[1635] = ~window[24][3];
assign temp[1636] = ~window[24][4];
assign temp[1637] = ~window[24][5];
assign temp[1638] = ~window[24][6];
assign temp[1639] = window[24][7];
assign temp[1640] = ~window[24][8];
assign temp[1664] = ~window[25][0];
assign temp[1665] = ~window[25][1];
assign temp[1666] = ~window[25][2];
assign temp[1667] = window[25][3];
assign temp[1668] = window[25][4];
assign temp[1669] = ~window[25][5];
assign temp[1670] = ~window[25][6];
assign temp[1671] = window[25][7];
assign temp[1672] = ~window[25][8];
assign temp[1696] = window[26][0];
assign temp[1697] = window[26][1];
assign temp[1698] = window[26][2];
assign temp[1699] = window[26][3];
assign temp[1700] = ~window[26][4];
assign temp[1701] = window[26][5];
assign temp[1702] = window[26][6];
assign temp[1703] = ~window[26][7];
assign temp[1704] = window[26][8];
assign temp[1728] = window[27][0];
assign temp[1729] = window[27][1];
assign temp[1730] = ~window[27][2];
assign temp[1731] = ~window[27][3];
assign temp[1732] = window[27][4];
assign temp[1733] = window[27][5];
assign temp[1734] = ~window[27][6];
assign temp[1735] = window[27][7];
assign temp[1736] = window[27][8];
assign temp[1760] = window[28][0];
assign temp[1761] = window[28][1];
assign temp[1762] = ~window[28][2];
assign temp[1763] = ~window[28][3];
assign temp[1764] = window[28][4];
assign temp[1765] = window[28][5];
assign temp[1766] = ~window[28][6];
assign temp[1767] = ~window[28][7];
assign temp[1768] = ~window[28][8];
assign temp[1792] = window[29][0];
assign temp[1793] = window[29][1];
assign temp[1794] = ~window[29][2];
assign temp[1795] = ~window[29][3];
assign temp[1796] = window[29][4];
assign temp[1797] = ~window[29][5];
assign temp[1798] = ~window[29][6];
assign temp[1799] = ~window[29][7];
assign temp[1800] = window[29][8];
assign temp[1824] = ~window[30][0];
assign temp[1825] = ~window[30][1];
assign temp[1826] = ~window[30][2];
assign temp[1827] = ~window[30][3];
assign temp[1828] = ~window[30][4];
assign temp[1829] = ~window[30][5];
assign temp[1830] = ~window[30][6];
assign temp[1831] = ~window[30][7];
assign temp[1832] = ~window[30][8];
assign temp[1856] = ~window[31][0];
assign temp[1857] = ~window[31][1];
assign temp[1858] = ~window[31][2];
assign temp[1859] = ~window[31][3];
assign temp[1860] = ~window[31][4];
assign temp[1861] = ~window[31][5];
assign temp[1862] = ~window[31][6];
assign temp[1863] = ~window[31][7];
assign temp[1864] = ~window[31][8];
assign temp[896] = ~window[0][0];
assign temp[897] = window[0][1];
assign temp[898] = window[0][2];
assign temp[899] = ~window[0][3];
assign temp[900] = ~window[0][4];
assign temp[901] = ~window[0][5];
assign temp[902] = window[0][6];
assign temp[903] = window[0][7];
assign temp[904] = window[0][8];
assign temp[928] = ~window[1][0];
assign temp[929] = ~window[1][1];
assign temp[930] = ~window[1][2];
assign temp[931] = ~window[1][3];
assign temp[932] = ~window[1][4];
assign temp[933] = ~window[1][5];
assign temp[934] = window[1][6];
assign temp[935] = window[1][7];
assign temp[936] = window[1][8];
assign temp[960] = window[2][0];
assign temp[961] = window[2][1];
assign temp[962] = window[2][2];
assign temp[963] = ~window[2][3];
assign temp[964] = window[2][4];
assign temp[965] = window[2][5];
assign temp[966] = ~window[2][6];
assign temp[967] = ~window[2][7];
assign temp[968] = ~window[2][8];
assign temp[992] = ~window[3][0];
assign temp[993] = ~window[3][1];
assign temp[994] = ~window[3][2];
assign temp[995] = ~window[3][3];
assign temp[996] = ~window[3][4];
assign temp[997] = ~window[3][5];
assign temp[998] = ~window[3][6];
assign temp[999] = window[3][7];
assign temp[1000] = window[3][8];
assign temp[1024] = window[4][0];
assign temp[1025] = ~window[4][1];
assign temp[1026] = window[4][2];
assign temp[1027] = window[4][3];
assign temp[1028] = window[4][4];
assign temp[1029] = window[4][5];
assign temp[1030] = ~window[4][6];
assign temp[1031] = ~window[4][7];
assign temp[1032] = window[4][8];
assign temp[1056] = ~window[5][0];
assign temp[1057] = ~window[5][1];
assign temp[1058] = ~window[5][2];
assign temp[1059] = window[5][3];
assign temp[1060] = ~window[5][4];
assign temp[1061] = ~window[5][5];
assign temp[1062] = window[5][6];
assign temp[1063] = ~window[5][7];
assign temp[1064] = window[5][8];
assign temp[1088] = window[6][0];
assign temp[1089] = window[6][1];
assign temp[1090] = window[6][2];
assign temp[1091] = window[6][3];
assign temp[1092] = ~window[6][4];
assign temp[1093] = window[6][5];
assign temp[1094] = ~window[6][6];
assign temp[1095] = ~window[6][7];
assign temp[1096] = window[6][8];
assign temp[1120] = ~window[7][0];
assign temp[1121] = ~window[7][1];
assign temp[1122] = ~window[7][2];
assign temp[1123] = window[7][3];
assign temp[1124] = window[7][4];
assign temp[1125] = window[7][5];
assign temp[1126] = window[7][6];
assign temp[1127] = ~window[7][7];
assign temp[1128] = ~window[7][8];
assign temp[1152] = window[8][0];
assign temp[1153] = window[8][1];
assign temp[1154] = window[8][2];
assign temp[1155] = window[8][3];
assign temp[1156] = window[8][4];
assign temp[1157] = ~window[8][5];
assign temp[1158] = window[8][6];
assign temp[1159] = window[8][7];
assign temp[1160] = window[8][8];
assign temp[1184] = ~window[9][0];
assign temp[1185] = ~window[9][1];
assign temp[1186] = ~window[9][2];
assign temp[1187] = ~window[9][3];
assign temp[1188] = ~window[9][4];
assign temp[1189] = ~window[9][5];
assign temp[1190] = window[9][6];
assign temp[1191] = window[9][7];
assign temp[1192] = window[9][8];
assign temp[1216] = ~window[10][0];
assign temp[1217] = ~window[10][1];
assign temp[1218] = ~window[10][2];
assign temp[1219] = window[10][3];
assign temp[1220] = window[10][4];
assign temp[1221] = ~window[10][5];
assign temp[1222] = ~window[10][6];
assign temp[1223] = ~window[10][7];
assign temp[1224] = window[10][8];
assign temp[1248] = window[11][0];
assign temp[1249] = window[11][1];
assign temp[1250] = window[11][2];
assign temp[1251] = window[11][3];
assign temp[1252] = ~window[11][4];
assign temp[1253] = window[11][5];
assign temp[1254] = window[11][6];
assign temp[1255] = ~window[11][7];
assign temp[1256] = ~window[11][8];
assign temp[1280] = window[12][0];
assign temp[1281] = window[12][1];
assign temp[1282] = window[12][2];
assign temp[1283] = window[12][3];
assign temp[1284] = ~window[12][4];
assign temp[1285] = window[12][5];
assign temp[1286] = ~window[12][6];
assign temp[1287] = ~window[12][7];
assign temp[1288] = ~window[12][8];
assign temp[1312] = ~window[13][0];
assign temp[1313] = ~window[13][1];
assign temp[1314] = ~window[13][2];
assign temp[1315] = window[13][3];
assign temp[1316] = ~window[13][4];
assign temp[1317] = ~window[13][5];
assign temp[1318] = window[13][6];
assign temp[1319] = window[13][7];
assign temp[1320] = ~window[13][8];
assign temp[1344] = ~window[14][0];
assign temp[1345] = ~window[14][1];
assign temp[1346] = ~window[14][2];
assign temp[1347] = window[14][3];
assign temp[1348] = ~window[14][4];
assign temp[1349] = ~window[14][5];
assign temp[1350] = ~window[14][6];
assign temp[1351] = window[14][7];
assign temp[1352] = window[14][8];
assign temp[1376] = ~window[15][0];
assign temp[1377] = ~window[15][1];
assign temp[1378] = ~window[15][2];
assign temp[1379] = ~window[15][3];
assign temp[1380] = window[15][4];
assign temp[1381] = ~window[15][5];
assign temp[1382] = ~window[15][6];
assign temp[1383] = ~window[15][7];
assign temp[1384] = ~window[15][8];
assign temp[1408] = ~window[16][0];
assign temp[1409] = ~window[16][1];
assign temp[1410] = ~window[16][2];
assign temp[1411] = ~window[16][3];
assign temp[1412] = window[16][4];
assign temp[1413] = window[16][5];
assign temp[1414] = ~window[16][6];
assign temp[1415] = ~window[16][7];
assign temp[1416] = ~window[16][8];
assign temp[1440] = ~window[17][0];
assign temp[1441] = ~window[17][1];
assign temp[1442] = window[17][2];
assign temp[1443] = window[17][3];
assign temp[1444] = ~window[17][4];
assign temp[1445] = ~window[17][5];
assign temp[1446] = window[17][6];
assign temp[1447] = window[17][7];
assign temp[1448] = window[17][8];
assign temp[1472] = ~window[18][0];
assign temp[1473] = window[18][1];
assign temp[1474] = ~window[18][2];
assign temp[1475] = window[18][3];
assign temp[1476] = window[18][4];
assign temp[1477] = ~window[18][5];
assign temp[1478] = ~window[18][6];
assign temp[1479] = window[18][7];
assign temp[1480] = window[18][8];
assign temp[1504] = ~window[19][0];
assign temp[1505] = ~window[19][1];
assign temp[1506] = window[19][2];
assign temp[1507] = window[19][3];
assign temp[1508] = ~window[19][4];
assign temp[1509] = ~window[19][5];
assign temp[1510] = window[19][6];
assign temp[1511] = window[19][7];
assign temp[1512] = ~window[19][8];
assign temp[1536] = ~window[20][0];
assign temp[1537] = ~window[20][1];
assign temp[1538] = ~window[20][2];
assign temp[1539] = ~window[20][3];
assign temp[1540] = ~window[20][4];
assign temp[1541] = ~window[20][5];
assign temp[1542] = window[20][6];
assign temp[1543] = window[20][7];
assign temp[1544] = window[20][8];
assign temp[1568] = ~window[21][0];
assign temp[1569] = ~window[21][1];
assign temp[1570] = ~window[21][2];
assign temp[1571] = ~window[21][3];
assign temp[1572] = ~window[21][4];
assign temp[1573] = ~window[21][5];
assign temp[1574] = window[21][6];
assign temp[1575] = ~window[21][7];
assign temp[1576] = ~window[21][8];
assign temp[1600] = window[22][0];
assign temp[1601] = ~window[22][1];
assign temp[1602] = window[22][2];
assign temp[1603] = window[22][3];
assign temp[1604] = window[22][4];
assign temp[1605] = window[22][5];
assign temp[1606] = ~window[22][6];
assign temp[1607] = ~window[22][7];
assign temp[1608] = ~window[22][8];
assign temp[1632] = ~window[23][0];
assign temp[1633] = ~window[23][1];
assign temp[1634] = ~window[23][2];
assign temp[1635] = ~window[23][3];
assign temp[1636] = ~window[23][4];
assign temp[1637] = ~window[23][5];
assign temp[1638] = window[23][6];
assign temp[1639] = window[23][7];
assign temp[1640] = window[23][8];
assign temp[1664] = window[24][0];
assign temp[1665] = window[24][1];
assign temp[1666] = window[24][2];
assign temp[1667] = ~window[24][3];
assign temp[1668] = ~window[24][4];
assign temp[1669] = ~window[24][5];
assign temp[1670] = ~window[24][6];
assign temp[1671] = window[24][7];
assign temp[1672] = window[24][8];
assign temp[1696] = ~window[25][0];
assign temp[1697] = ~window[25][1];
assign temp[1698] = ~window[25][2];
assign temp[1699] = ~window[25][3];
assign temp[1700] = window[25][4];
assign temp[1701] = ~window[25][5];
assign temp[1702] = window[25][6];
assign temp[1703] = window[25][7];
assign temp[1704] = ~window[25][8];
assign temp[1728] = ~window[26][0];
assign temp[1729] = window[26][1];
assign temp[1730] = window[26][2];
assign temp[1731] = ~window[26][3];
assign temp[1732] = ~window[26][4];
assign temp[1733] = ~window[26][5];
assign temp[1734] = window[26][6];
assign temp[1735] = ~window[26][7];
assign temp[1736] = ~window[26][8];
assign temp[1760] = ~window[27][0];
assign temp[1761] = ~window[27][1];
assign temp[1762] = window[27][2];
assign temp[1763] = window[27][3];
assign temp[1764] = window[27][4];
assign temp[1765] = window[27][5];
assign temp[1766] = ~window[27][6];
assign temp[1767] = ~window[27][7];
assign temp[1768] = ~window[27][8];
assign temp[1792] = window[28][0];
assign temp[1793] = window[28][1];
assign temp[1794] = ~window[28][2];
assign temp[1795] = window[28][3];
assign temp[1796] = ~window[28][4];
assign temp[1797] = ~window[28][5];
assign temp[1798] = ~window[28][6];
assign temp[1799] = ~window[28][7];
assign temp[1800] = ~window[28][8];
assign temp[1824] = window[29][0];
assign temp[1825] = ~window[29][1];
assign temp[1826] = window[29][2];
assign temp[1827] = window[29][3];
assign temp[1828] = window[29][4];
assign temp[1829] = window[29][5];
assign temp[1830] = ~window[29][6];
assign temp[1831] = window[29][7];
assign temp[1832] = window[29][8];
assign temp[1856] = ~window[30][0];
assign temp[1857] = ~window[30][1];
assign temp[1858] = ~window[30][2];
assign temp[1859] = window[30][3];
assign temp[1860] = ~window[30][4];
assign temp[1861] = window[30][5];
assign temp[1862] = ~window[30][6];
assign temp[1863] = window[30][7];
assign temp[1864] = window[30][8];
assign temp[1888] = window[31][0];
assign temp[1889] = window[31][1];
assign temp[1890] = window[31][2];
assign temp[1891] = window[31][3];
assign temp[1892] = ~window[31][4];
assign temp[1893] = ~window[31][5];
assign temp[1894] = window[31][6];
assign temp[1895] = ~window[31][7];
assign temp[1896] = ~window[31][8];
assign temp[928] = ~window[0][0];
assign temp[929] = ~window[0][1];
assign temp[930] = window[0][2];
assign temp[931] = window[0][3];
assign temp[932] = window[0][4];
assign temp[933] = window[0][5];
assign temp[934] = ~window[0][6];
assign temp[935] = ~window[0][7];
assign temp[936] = window[0][8];
assign temp[960] = ~window[1][0];
assign temp[961] = ~window[1][1];
assign temp[962] = window[1][2];
assign temp[963] = window[1][3];
assign temp[964] = window[1][4];
assign temp[965] = window[1][5];
assign temp[966] = ~window[1][6];
assign temp[967] = ~window[1][7];
assign temp[968] = window[1][8];
assign temp[992] = window[2][0];
assign temp[993] = window[2][1];
assign temp[994] = window[2][2];
assign temp[995] = window[2][3];
assign temp[996] = window[2][4];
assign temp[997] = window[2][5];
assign temp[998] = window[2][6];
assign temp[999] = window[2][7];
assign temp[1000] = ~window[2][8];
assign temp[1024] = ~window[3][0];
assign temp[1025] = ~window[3][1];
assign temp[1026] = ~window[3][2];
assign temp[1027] = window[3][3];
assign temp[1028] = ~window[3][4];
assign temp[1029] = ~window[3][5];
assign temp[1030] = ~window[3][6];
assign temp[1031] = ~window[3][7];
assign temp[1032] = ~window[3][8];
assign temp[1056] = ~window[4][0];
assign temp[1057] = window[4][1];
assign temp[1058] = window[4][2];
assign temp[1059] = window[4][3];
assign temp[1060] = window[4][4];
assign temp[1061] = window[4][5];
assign temp[1062] = window[4][6];
assign temp[1063] = window[4][7];
assign temp[1064] = window[4][8];
assign temp[1088] = ~window[5][0];
assign temp[1089] = window[5][1];
assign temp[1090] = ~window[5][2];
assign temp[1091] = window[5][3];
assign temp[1092] = window[5][4];
assign temp[1093] = ~window[5][5];
assign temp[1094] = ~window[5][6];
assign temp[1095] = window[5][7];
assign temp[1096] = window[5][8];
assign temp[1120] = window[6][0];
assign temp[1121] = ~window[6][1];
assign temp[1122] = window[6][2];
assign temp[1123] = window[6][3];
assign temp[1124] = window[6][4];
assign temp[1125] = window[6][5];
assign temp[1126] = window[6][6];
assign temp[1127] = window[6][7];
assign temp[1128] = window[6][8];
assign temp[1152] = ~window[7][0];
assign temp[1153] = ~window[7][1];
assign temp[1154] = ~window[7][2];
assign temp[1155] = ~window[7][3];
assign temp[1156] = window[7][4];
assign temp[1157] = ~window[7][5];
assign temp[1158] = window[7][6];
assign temp[1159] = window[7][7];
assign temp[1160] = ~window[7][8];
assign temp[1184] = ~window[8][0];
assign temp[1185] = window[8][1];
assign temp[1186] = ~window[8][2];
assign temp[1187] = window[8][3];
assign temp[1188] = window[8][4];
assign temp[1189] = window[8][5];
assign temp[1190] = ~window[8][6];
assign temp[1191] = ~window[8][7];
assign temp[1192] = ~window[8][8];
assign temp[1216] = window[9][0];
assign temp[1217] = window[9][1];
assign temp[1218] = window[9][2];
assign temp[1219] = ~window[9][3];
assign temp[1220] = ~window[9][4];
assign temp[1221] = ~window[9][5];
assign temp[1222] = ~window[9][6];
assign temp[1223] = ~window[9][7];
assign temp[1224] = ~window[9][8];
assign temp[1248] = ~window[10][0];
assign temp[1249] = ~window[10][1];
assign temp[1250] = ~window[10][2];
assign temp[1251] = ~window[10][3];
assign temp[1252] = ~window[10][4];
assign temp[1253] = window[10][5];
assign temp[1254] = window[10][6];
assign temp[1255] = window[10][7];
assign temp[1256] = window[10][8];
assign temp[1280] = window[11][0];
assign temp[1281] = window[11][1];
assign temp[1282] = window[11][2];
assign temp[1283] = window[11][3];
assign temp[1284] = window[11][4];
assign temp[1285] = window[11][5];
assign temp[1286] = window[11][6];
assign temp[1287] = ~window[11][7];
assign temp[1288] = window[11][8];
assign temp[1312] = window[12][0];
assign temp[1313] = ~window[12][1];
assign temp[1314] = ~window[12][2];
assign temp[1315] = window[12][3];
assign temp[1316] = window[12][4];
assign temp[1317] = window[12][5];
assign temp[1318] = window[12][6];
assign temp[1319] = ~window[12][7];
assign temp[1320] = ~window[12][8];
assign temp[1344] = ~window[13][0];
assign temp[1345] = ~window[13][1];
assign temp[1346] = ~window[13][2];
assign temp[1347] = ~window[13][3];
assign temp[1348] = window[13][4];
assign temp[1349] = ~window[13][5];
assign temp[1350] = ~window[13][6];
assign temp[1351] = ~window[13][7];
assign temp[1352] = ~window[13][8];
assign temp[1376] = ~window[14][0];
assign temp[1377] = ~window[14][1];
assign temp[1378] = ~window[14][2];
assign temp[1379] = window[14][3];
assign temp[1380] = window[14][4];
assign temp[1381] = window[14][5];
assign temp[1382] = ~window[14][6];
assign temp[1383] = ~window[14][7];
assign temp[1384] = ~window[14][8];
assign temp[1408] = window[15][0];
assign temp[1409] = window[15][1];
assign temp[1410] = window[15][2];
assign temp[1411] = window[15][3];
assign temp[1412] = ~window[15][4];
assign temp[1413] = window[15][5];
assign temp[1414] = window[15][6];
assign temp[1415] = window[15][7];
assign temp[1416] = window[15][8];
assign temp[1440] = ~window[16][0];
assign temp[1441] = window[16][1];
assign temp[1442] = ~window[16][2];
assign temp[1443] = window[16][3];
assign temp[1444] = window[16][4];
assign temp[1445] = ~window[16][5];
assign temp[1446] = ~window[16][6];
assign temp[1447] = ~window[16][7];
assign temp[1448] = ~window[16][8];
assign temp[1472] = ~window[17][0];
assign temp[1473] = window[17][1];
assign temp[1474] = window[17][2];
assign temp[1475] = window[17][3];
assign temp[1476] = window[17][4];
assign temp[1477] = window[17][5];
assign temp[1478] = ~window[17][6];
assign temp[1479] = window[17][7];
assign temp[1480] = ~window[17][8];
assign temp[1504] = window[18][0];
assign temp[1505] = window[18][1];
assign temp[1506] = window[18][2];
assign temp[1507] = ~window[18][3];
assign temp[1508] = ~window[18][4];
assign temp[1509] = ~window[18][5];
assign temp[1510] = window[18][6];
assign temp[1511] = window[18][7];
assign temp[1512] = window[18][8];
assign temp[1536] = ~window[19][0];
assign temp[1537] = window[19][1];
assign temp[1538] = window[19][2];
assign temp[1539] = window[19][3];
assign temp[1540] = ~window[19][4];
assign temp[1541] = window[19][5];
assign temp[1542] = window[19][6];
assign temp[1543] = window[19][7];
assign temp[1544] = window[19][8];
assign temp[1568] = ~window[20][0];
assign temp[1569] = ~window[20][1];
assign temp[1570] = ~window[20][2];
assign temp[1571] = ~window[20][3];
assign temp[1572] = ~window[20][4];
assign temp[1573] = ~window[20][5];
assign temp[1574] = ~window[20][6];
assign temp[1575] = ~window[20][7];
assign temp[1576] = ~window[20][8];
assign temp[1600] = ~window[21][0];
assign temp[1601] = ~window[21][1];
assign temp[1602] = ~window[21][2];
assign temp[1603] = window[21][3];
assign temp[1604] = ~window[21][4];
assign temp[1605] = window[21][5];
assign temp[1606] = window[21][6];
assign temp[1607] = window[21][7];
assign temp[1608] = ~window[21][8];
assign temp[1632] = window[22][0];
assign temp[1633] = window[22][1];
assign temp[1634] = ~window[22][2];
assign temp[1635] = window[22][3];
assign temp[1636] = window[22][4];
assign temp[1637] = window[22][5];
assign temp[1638] = window[22][6];
assign temp[1639] = window[22][7];
assign temp[1640] = window[22][8];
assign temp[1664] = ~window[23][0];
assign temp[1665] = window[23][1];
assign temp[1666] = ~window[23][2];
assign temp[1667] = ~window[23][3];
assign temp[1668] = window[23][4];
assign temp[1669] = ~window[23][5];
assign temp[1670] = ~window[23][6];
assign temp[1671] = ~window[23][7];
assign temp[1672] = ~window[23][8];
assign temp[1696] = window[24][0];
assign temp[1697] = window[24][1];
assign temp[1698] = window[24][2];
assign temp[1699] = window[24][3];
assign temp[1700] = window[24][4];
assign temp[1701] = window[24][5];
assign temp[1702] = ~window[24][6];
assign temp[1703] = window[24][7];
assign temp[1704] = ~window[24][8];
assign temp[1728] = ~window[25][0];
assign temp[1729] = window[25][1];
assign temp[1730] = ~window[25][2];
assign temp[1731] = ~window[25][3];
assign temp[1732] = window[25][4];
assign temp[1733] = window[25][5];
assign temp[1734] = window[25][6];
assign temp[1735] = ~window[25][7];
assign temp[1736] = ~window[25][8];
assign temp[1760] = ~window[26][0];
assign temp[1761] = ~window[26][1];
assign temp[1762] = window[26][2];
assign temp[1763] = window[26][3];
assign temp[1764] = window[26][4];
assign temp[1765] = window[26][5];
assign temp[1766] = window[26][6];
assign temp[1767] = window[26][7];
assign temp[1768] = window[26][8];
assign temp[1792] = ~window[27][0];
assign temp[1793] = ~window[27][1];
assign temp[1794] = window[27][2];
assign temp[1795] = ~window[27][3];
assign temp[1796] = ~window[27][4];
assign temp[1797] = ~window[27][5];
assign temp[1798] = window[27][6];
assign temp[1799] = window[27][7];
assign temp[1800] = window[27][8];
assign temp[1824] = ~window[28][0];
assign temp[1825] = ~window[28][1];
assign temp[1826] = ~window[28][2];
assign temp[1827] = window[28][3];
assign temp[1828] = window[28][4];
assign temp[1829] = ~window[28][5];
assign temp[1830] = ~window[28][6];
assign temp[1831] = window[28][7];
assign temp[1832] = ~window[28][8];
assign temp[1856] = ~window[29][0];
assign temp[1857] = ~window[29][1];
assign temp[1858] = ~window[29][2];
assign temp[1859] = ~window[29][3];
assign temp[1860] = window[29][4];
assign temp[1861] = window[29][5];
assign temp[1862] = ~window[29][6];
assign temp[1863] = ~window[29][7];
assign temp[1864] = ~window[29][8];
assign temp[1888] = ~window[30][0];
assign temp[1889] = window[30][1];
assign temp[1890] = ~window[30][2];
assign temp[1891] = ~window[30][3];
assign temp[1892] = window[30][4];
assign temp[1893] = ~window[30][5];
assign temp[1894] = ~window[30][6];
assign temp[1895] = window[30][7];
assign temp[1896] = window[30][8];
assign temp[1920] = window[31][0];
assign temp[1921] = window[31][1];
assign temp[1922] = window[31][2];
assign temp[1923] = window[31][3];
assign temp[1924] = window[31][4];
assign temp[1925] = window[31][5];
assign temp[1926] = ~window[31][6];
assign temp[1927] = window[31][7];
assign temp[1928] = ~window[31][8];
assign temp[960] = ~window[0][0];
assign temp[961] = ~window[0][1];
assign temp[962] = ~window[0][2];
assign temp[963] = ~window[0][3];
assign temp[964] = ~window[0][4];
assign temp[965] = ~window[0][5];
assign temp[966] = ~window[0][6];
assign temp[967] = ~window[0][7];
assign temp[968] = ~window[0][8];
assign temp[992] = window[1][0];
assign temp[993] = window[1][1];
assign temp[994] = window[1][2];
assign temp[995] = window[1][3];
assign temp[996] = window[1][4];
assign temp[997] = window[1][5];
assign temp[998] = window[1][6];
assign temp[999] = ~window[1][7];
assign temp[1000] = window[1][8];
assign temp[1024] = ~window[2][0];
assign temp[1025] = ~window[2][1];
assign temp[1026] = window[2][2];
assign temp[1027] = ~window[2][3];
assign temp[1028] = ~window[2][4];
assign temp[1029] = ~window[2][5];
assign temp[1030] = ~window[2][6];
assign temp[1031] = ~window[2][7];
assign temp[1032] = ~window[2][8];
assign temp[1056] = window[3][0];
assign temp[1057] = window[3][1];
assign temp[1058] = window[3][2];
assign temp[1059] = window[3][3];
assign temp[1060] = window[3][4];
assign temp[1061] = window[3][5];
assign temp[1062] = window[3][6];
assign temp[1063] = window[3][7];
assign temp[1064] = window[3][8];
assign temp[1088] = window[4][0];
assign temp[1089] = ~window[4][1];
assign temp[1090] = ~window[4][2];
assign temp[1091] = ~window[4][3];
assign temp[1092] = window[4][4];
assign temp[1093] = window[4][5];
assign temp[1094] = window[4][6];
assign temp[1095] = window[4][7];
assign temp[1096] = window[4][8];
assign temp[1120] = window[5][0];
assign temp[1121] = window[5][1];
assign temp[1122] = ~window[5][2];
assign temp[1123] = window[5][3];
assign temp[1124] = window[5][4];
assign temp[1125] = ~window[5][5];
assign temp[1126] = window[5][6];
assign temp[1127] = window[5][7];
assign temp[1128] = window[5][8];
assign temp[1152] = ~window[6][0];
assign temp[1153] = ~window[6][1];
assign temp[1154] = ~window[6][2];
assign temp[1155] = ~window[6][3];
assign temp[1156] = ~window[6][4];
assign temp[1157] = window[6][5];
assign temp[1158] = window[6][6];
assign temp[1159] = ~window[6][7];
assign temp[1160] = ~window[6][8];
assign temp[1184] = window[7][0];
assign temp[1185] = window[7][1];
assign temp[1186] = window[7][2];
assign temp[1187] = window[7][3];
assign temp[1188] = window[7][4];
assign temp[1189] = window[7][5];
assign temp[1190] = window[7][6];
assign temp[1191] = window[7][7];
assign temp[1192] = window[7][8];
assign temp[1216] = ~window[8][0];
assign temp[1217] = window[8][1];
assign temp[1218] = ~window[8][2];
assign temp[1219] = ~window[8][3];
assign temp[1220] = ~window[8][4];
assign temp[1221] = ~window[8][5];
assign temp[1222] = ~window[8][6];
assign temp[1223] = ~window[8][7];
assign temp[1224] = ~window[8][8];
assign temp[1248] = window[9][0];
assign temp[1249] = window[9][1];
assign temp[1250] = window[9][2];
assign temp[1251] = window[9][3];
assign temp[1252] = window[9][4];
assign temp[1253] = ~window[9][5];
assign temp[1254] = window[9][6];
assign temp[1255] = ~window[9][7];
assign temp[1256] = window[9][8];
assign temp[1280] = window[10][0];
assign temp[1281] = window[10][1];
assign temp[1282] = window[10][2];
assign temp[1283] = window[10][3];
assign temp[1284] = window[10][4];
assign temp[1285] = window[10][5];
assign temp[1286] = window[10][6];
assign temp[1287] = ~window[10][7];
assign temp[1288] = ~window[10][8];
assign temp[1312] = ~window[11][0];
assign temp[1313] = ~window[11][1];
assign temp[1314] = window[11][2];
assign temp[1315] = ~window[11][3];
assign temp[1316] = ~window[11][4];
assign temp[1317] = ~window[11][5];
assign temp[1318] = ~window[11][6];
assign temp[1319] = ~window[11][7];
assign temp[1320] = ~window[11][8];
assign temp[1344] = ~window[12][0];
assign temp[1345] = ~window[12][1];
assign temp[1346] = ~window[12][2];
assign temp[1347] = ~window[12][3];
assign temp[1348] = ~window[12][4];
assign temp[1349] = window[12][5];
assign temp[1350] = ~window[12][6];
assign temp[1351] = ~window[12][7];
assign temp[1352] = ~window[12][8];
assign temp[1376] = window[13][0];
assign temp[1377] = window[13][1];
assign temp[1378] = ~window[13][2];
assign temp[1379] = window[13][3];
assign temp[1380] = ~window[13][4];
assign temp[1381] = window[13][5];
assign temp[1382] = ~window[13][6];
assign temp[1383] = window[13][7];
assign temp[1384] = window[13][8];
assign temp[1408] = window[14][0];
assign temp[1409] = ~window[14][1];
assign temp[1410] = ~window[14][2];
assign temp[1411] = ~window[14][3];
assign temp[1412] = ~window[14][4];
assign temp[1413] = ~window[14][5];
assign temp[1414] = ~window[14][6];
assign temp[1415] = ~window[14][7];
assign temp[1416] = ~window[14][8];
assign temp[1440] = ~window[15][0];
assign temp[1441] = ~window[15][1];
assign temp[1442] = window[15][2];
assign temp[1443] = ~window[15][3];
assign temp[1444] = window[15][4];
assign temp[1445] = window[15][5];
assign temp[1446] = window[15][6];
assign temp[1447] = ~window[15][7];
assign temp[1448] = window[15][8];
assign temp[1472] = window[16][0];
assign temp[1473] = window[16][1];
assign temp[1474] = ~window[16][2];
assign temp[1475] = window[16][3];
assign temp[1476] = ~window[16][4];
assign temp[1477] = ~window[16][5];
assign temp[1478] = window[16][6];
assign temp[1479] = window[16][7];
assign temp[1480] = ~window[16][8];
assign temp[1504] = window[17][0];
assign temp[1505] = window[17][1];
assign temp[1506] = window[17][2];
assign temp[1507] = window[17][3];
assign temp[1508] = window[17][4];
assign temp[1509] = window[17][5];
assign temp[1510] = ~window[17][6];
assign temp[1511] = window[17][7];
assign temp[1512] = window[17][8];
assign temp[1536] = ~window[18][0];
assign temp[1537] = window[18][1];
assign temp[1538] = window[18][2];
assign temp[1539] = window[18][3];
assign temp[1540] = window[18][4];
assign temp[1541] = ~window[18][5];
assign temp[1542] = window[18][6];
assign temp[1543] = window[18][7];
assign temp[1544] = window[18][8];
assign temp[1568] = ~window[19][0];
assign temp[1569] = window[19][1];
assign temp[1570] = window[19][2];
assign temp[1571] = window[19][3];
assign temp[1572] = ~window[19][4];
assign temp[1573] = window[19][5];
assign temp[1574] = window[19][6];
assign temp[1575] = window[19][7];
assign temp[1576] = window[19][8];
assign temp[1600] = window[20][0];
assign temp[1601] = window[20][1];
assign temp[1602] = window[20][2];
assign temp[1603] = window[20][3];
assign temp[1604] = window[20][4];
assign temp[1605] = ~window[20][5];
assign temp[1606] = ~window[20][6];
assign temp[1607] = ~window[20][7];
assign temp[1608] = ~window[20][8];
assign temp[1632] = window[21][0];
assign temp[1633] = window[21][1];
assign temp[1634] = window[21][2];
assign temp[1635] = window[21][3];
assign temp[1636] = window[21][4];
assign temp[1637] = window[21][5];
assign temp[1638] = window[21][6];
assign temp[1639] = window[21][7];
assign temp[1640] = window[21][8];
assign temp[1664] = ~window[22][0];
assign temp[1665] = ~window[22][1];
assign temp[1666] = ~window[22][2];
assign temp[1667] = ~window[22][3];
assign temp[1668] = window[22][4];
assign temp[1669] = window[22][5];
assign temp[1670] = window[22][6];
assign temp[1671] = ~window[22][7];
assign temp[1672] = window[22][8];
assign temp[1696] = window[23][0];
assign temp[1697] = ~window[23][1];
assign temp[1698] = window[23][2];
assign temp[1699] = window[23][3];
assign temp[1700] = window[23][4];
assign temp[1701] = ~window[23][5];
assign temp[1702] = window[23][6];
assign temp[1703] = window[23][7];
assign temp[1704] = window[23][8];
assign temp[1728] = ~window[24][0];
assign temp[1729] = ~window[24][1];
assign temp[1730] = window[24][2];
assign temp[1731] = ~window[24][3];
assign temp[1732] = ~window[24][4];
assign temp[1733] = ~window[24][5];
assign temp[1734] = ~window[24][6];
assign temp[1735] = ~window[24][7];
assign temp[1736] = ~window[24][8];
assign temp[1760] = window[25][0];
assign temp[1761] = window[25][1];
assign temp[1762] = ~window[25][2];
assign temp[1763] = window[25][3];
assign temp[1764] = window[25][4];
assign temp[1765] = ~window[25][5];
assign temp[1766] = ~window[25][6];
assign temp[1767] = window[25][7];
assign temp[1768] = ~window[25][8];
assign temp[1792] = window[26][0];
assign temp[1793] = window[26][1];
assign temp[1794] = window[26][2];
assign temp[1795] = window[26][3];
assign temp[1796] = ~window[26][4];
assign temp[1797] = window[26][5];
assign temp[1798] = ~window[26][6];
assign temp[1799] = ~window[26][7];
assign temp[1800] = window[26][8];
assign temp[1824] = window[27][0];
assign temp[1825] = window[27][1];
assign temp[1826] = ~window[27][2];
assign temp[1827] = window[27][3];
assign temp[1828] = window[27][4];
assign temp[1829] = window[27][5];
assign temp[1830] = window[27][6];
assign temp[1831] = window[27][7];
assign temp[1832] = window[27][8];
assign temp[1856] = window[28][0];
assign temp[1857] = ~window[28][1];
assign temp[1858] = ~window[28][2];
assign temp[1859] = ~window[28][3];
assign temp[1860] = ~window[28][4];
assign temp[1861] = ~window[28][5];
assign temp[1862] = window[28][6];
assign temp[1863] = ~window[28][7];
assign temp[1864] = ~window[28][8];
assign temp[1888] = ~window[29][0];
assign temp[1889] = window[29][1];
assign temp[1890] = window[29][2];
assign temp[1891] = window[29][3];
assign temp[1892] = window[29][4];
assign temp[1893] = window[29][5];
assign temp[1894] = window[29][6];
assign temp[1895] = ~window[29][7];
assign temp[1896] = window[29][8];
assign temp[1920] = window[30][0];
assign temp[1921] = window[30][1];
assign temp[1922] = ~window[30][2];
assign temp[1923] = window[30][3];
assign temp[1924] = window[30][4];
assign temp[1925] = ~window[30][5];
assign temp[1926] = ~window[30][6];
assign temp[1927] = window[30][7];
assign temp[1928] = ~window[30][8];
assign temp[1952] = ~window[31][0];
assign temp[1953] = ~window[31][1];
assign temp[1954] = window[31][2];
assign temp[1955] = ~window[31][3];
assign temp[1956] = ~window[31][4];
assign temp[1957] = ~window[31][5];
assign temp[1958] = ~window[31][6];
assign temp[1959] = ~window[31][7];
assign temp[1960] = ~window[31][8];
assign temp[992] = window[0][0];
assign temp[993] = window[0][1];
assign temp[994] = ~window[0][2];
assign temp[995] = ~window[0][3];
assign temp[996] = ~window[0][4];
assign temp[997] = ~window[0][5];
assign temp[998] = ~window[0][6];
assign temp[999] = window[0][7];
assign temp[1000] = ~window[0][8];
assign temp[1024] = ~window[1][0];
assign temp[1025] = ~window[1][1];
assign temp[1026] = ~window[1][2];
assign temp[1027] = window[1][3];
assign temp[1028] = window[1][4];
assign temp[1029] = window[1][5];
assign temp[1030] = ~window[1][6];
assign temp[1031] = window[1][7];
assign temp[1032] = ~window[1][8];
assign temp[1056] = ~window[2][0];
assign temp[1057] = ~window[2][1];
assign temp[1058] = window[2][2];
assign temp[1059] = window[2][3];
assign temp[1060] = ~window[2][4];
assign temp[1061] = ~window[2][5];
assign temp[1062] = window[2][6];
assign temp[1063] = window[2][7];
assign temp[1064] = ~window[2][8];
assign temp[1088] = window[3][0];
assign temp[1089] = window[3][1];
assign temp[1090] = window[3][2];
assign temp[1091] = window[3][3];
assign temp[1092] = window[3][4];
assign temp[1093] = window[3][5];
assign temp[1094] = ~window[3][6];
assign temp[1095] = ~window[3][7];
assign temp[1096] = ~window[3][8];
assign temp[1120] = window[4][0];
assign temp[1121] = ~window[4][1];
assign temp[1122] = ~window[4][2];
assign temp[1123] = ~window[4][3];
assign temp[1124] = ~window[4][4];
assign temp[1125] = ~window[4][5];
assign temp[1126] = ~window[4][6];
assign temp[1127] = ~window[4][7];
assign temp[1128] = ~window[4][8];
assign temp[1152] = window[5][0];
assign temp[1153] = window[5][1];
assign temp[1154] = ~window[5][2];
assign temp[1155] = ~window[5][3];
assign temp[1156] = ~window[5][4];
assign temp[1157] = ~window[5][5];
assign temp[1158] = ~window[5][6];
assign temp[1159] = ~window[5][7];
assign temp[1160] = ~window[5][8];
assign temp[1184] = ~window[6][0];
assign temp[1185] = ~window[6][1];
assign temp[1186] = ~window[6][2];
assign temp[1187] = ~window[6][3];
assign temp[1188] = ~window[6][4];
assign temp[1189] = window[6][5];
assign temp[1190] = window[6][6];
assign temp[1191] = window[6][7];
assign temp[1192] = ~window[6][8];
assign temp[1216] = window[7][0];
assign temp[1217] = window[7][1];
assign temp[1218] = window[7][2];
assign temp[1219] = ~window[7][3];
assign temp[1220] = ~window[7][4];
assign temp[1221] = ~window[7][5];
assign temp[1222] = ~window[7][6];
assign temp[1223] = ~window[7][7];
assign temp[1224] = ~window[7][8];
assign temp[1248] = window[8][0];
assign temp[1249] = ~window[8][1];
assign temp[1250] = ~window[8][2];
assign temp[1251] = ~window[8][3];
assign temp[1252] = ~window[8][4];
assign temp[1253] = ~window[8][5];
assign temp[1254] = ~window[8][6];
assign temp[1255] = ~window[8][7];
assign temp[1256] = ~window[8][8];
assign temp[1280] = window[9][0];
assign temp[1281] = window[9][1];
assign temp[1282] = window[9][2];
assign temp[1283] = window[9][3];
assign temp[1284] = window[9][4];
assign temp[1285] = ~window[9][5];
assign temp[1286] = ~window[9][6];
assign temp[1287] = window[9][7];
assign temp[1288] = ~window[9][8];
assign temp[1312] = window[10][0];
assign temp[1313] = window[10][1];
assign temp[1314] = window[10][2];
assign temp[1315] = window[10][3];
assign temp[1316] = window[10][4];
assign temp[1317] = window[10][5];
assign temp[1318] = ~window[10][6];
assign temp[1319] = ~window[10][7];
assign temp[1320] = ~window[10][8];
assign temp[1344] = window[11][0];
assign temp[1345] = window[11][1];
assign temp[1346] = ~window[11][2];
assign temp[1347] = window[11][3];
assign temp[1348] = ~window[11][4];
assign temp[1349] = ~window[11][5];
assign temp[1350] = ~window[11][6];
assign temp[1351] = window[11][7];
assign temp[1352] = window[11][8];
assign temp[1376] = ~window[12][0];
assign temp[1377] = ~window[12][1];
assign temp[1378] = window[12][2];
assign temp[1379] = window[12][3];
assign temp[1380] = ~window[12][4];
assign temp[1381] = window[12][5];
assign temp[1382] = window[12][6];
assign temp[1383] = window[12][7];
assign temp[1384] = window[12][8];
assign temp[1408] = ~window[13][0];
assign temp[1409] = window[13][1];
assign temp[1410] = window[13][2];
assign temp[1411] = ~window[13][3];
assign temp[1412] = window[13][4];
assign temp[1413] = window[13][5];
assign temp[1414] = ~window[13][6];
assign temp[1415] = window[13][7];
assign temp[1416] = window[13][8];
assign temp[1440] = window[14][0];
assign temp[1441] = window[14][1];
assign temp[1442] = ~window[14][2];
assign temp[1443] = ~window[14][3];
assign temp[1444] = ~window[14][4];
assign temp[1445] = ~window[14][5];
assign temp[1446] = ~window[14][6];
assign temp[1447] = ~window[14][7];
assign temp[1448] = window[14][8];
assign temp[1472] = ~window[15][0];
assign temp[1473] = ~window[15][1];
assign temp[1474] = ~window[15][2];
assign temp[1475] = ~window[15][3];
assign temp[1476] = ~window[15][4];
assign temp[1477] = ~window[15][5];
assign temp[1478] = ~window[15][6];
assign temp[1479] = window[15][7];
assign temp[1480] = window[15][8];
assign temp[1504] = ~window[16][0];
assign temp[1505] = ~window[16][1];
assign temp[1506] = ~window[16][2];
assign temp[1507] = ~window[16][3];
assign temp[1508] = ~window[16][4];
assign temp[1509] = ~window[16][5];
assign temp[1510] = ~window[16][6];
assign temp[1511] = ~window[16][7];
assign temp[1512] = window[16][8];
assign temp[1536] = ~window[17][0];
assign temp[1537] = ~window[17][1];
assign temp[1538] = window[17][2];
assign temp[1539] = window[17][3];
assign temp[1540] = window[17][4];
assign temp[1541] = window[17][5];
assign temp[1542] = window[17][6];
assign temp[1543] = window[17][7];
assign temp[1544] = ~window[17][8];
assign temp[1568] = ~window[18][0];
assign temp[1569] = ~window[18][1];
assign temp[1570] = window[18][2];
assign temp[1571] = ~window[18][3];
assign temp[1572] = ~window[18][4];
assign temp[1573] = ~window[18][5];
assign temp[1574] = ~window[18][6];
assign temp[1575] = ~window[18][7];
assign temp[1576] = window[18][8];
assign temp[1600] = window[19][0];
assign temp[1601] = ~window[19][1];
assign temp[1602] = ~window[19][2];
assign temp[1603] = window[19][3];
assign temp[1604] = window[19][4];
assign temp[1605] = window[19][5];
assign temp[1606] = ~window[19][6];
assign temp[1607] = window[19][7];
assign temp[1608] = window[19][8];
assign temp[1632] = ~window[20][0];
assign temp[1633] = window[20][1];
assign temp[1634] = window[20][2];
assign temp[1635] = window[20][3];
assign temp[1636] = window[20][4];
assign temp[1637] = ~window[20][5];
assign temp[1638] = window[20][6];
assign temp[1639] = ~window[20][7];
assign temp[1640] = ~window[20][8];
assign temp[1664] = ~window[21][0];
assign temp[1665] = window[21][1];
assign temp[1666] = ~window[21][2];
assign temp[1667] = window[21][3];
assign temp[1668] = window[21][4];
assign temp[1669] = window[21][5];
assign temp[1670] = ~window[21][6];
assign temp[1671] = window[21][7];
assign temp[1672] = window[21][8];
assign temp[1696] = ~window[22][0];
assign temp[1697] = window[22][1];
assign temp[1698] = window[22][2];
assign temp[1699] = ~window[22][3];
assign temp[1700] = ~window[22][4];
assign temp[1701] = ~window[22][5];
assign temp[1702] = ~window[22][6];
assign temp[1703] = window[22][7];
assign temp[1704] = window[22][8];
assign temp[1728] = window[23][0];
assign temp[1729] = window[23][1];
assign temp[1730] = window[23][2];
assign temp[1731] = window[23][3];
assign temp[1732] = ~window[23][4];
assign temp[1733] = ~window[23][5];
assign temp[1734] = ~window[23][6];
assign temp[1735] = ~window[23][7];
assign temp[1736] = ~window[23][8];
assign temp[1760] = ~window[24][0];
assign temp[1761] = ~window[24][1];
assign temp[1762] = ~window[24][2];
assign temp[1763] = window[24][3];
assign temp[1764] = window[24][4];
assign temp[1765] = window[24][5];
assign temp[1766] = window[24][6];
assign temp[1767] = window[24][7];
assign temp[1768] = ~window[24][8];
assign temp[1792] = ~window[25][0];
assign temp[1793] = window[25][1];
assign temp[1794] = window[25][2];
assign temp[1795] = ~window[25][3];
assign temp[1796] = window[25][4];
assign temp[1797] = ~window[25][5];
assign temp[1798] = ~window[25][6];
assign temp[1799] = ~window[25][7];
assign temp[1800] = window[25][8];
assign temp[1824] = window[26][0];
assign temp[1825] = window[26][1];
assign temp[1826] = ~window[26][2];
assign temp[1827] = window[26][3];
assign temp[1828] = ~window[26][4];
assign temp[1829] = window[26][5];
assign temp[1830] = window[26][6];
assign temp[1831] = window[26][7];
assign temp[1832] = window[26][8];
assign temp[1856] = window[27][0];
assign temp[1857] = window[27][1];
assign temp[1858] = window[27][2];
assign temp[1859] = ~window[27][3];
assign temp[1860] = ~window[27][4];
assign temp[1861] = ~window[27][5];
assign temp[1862] = ~window[27][6];
assign temp[1863] = ~window[27][7];
assign temp[1864] = window[27][8];
assign temp[1888] = ~window[28][0];
assign temp[1889] = ~window[28][1];
assign temp[1890] = ~window[28][2];
assign temp[1891] = ~window[28][3];
assign temp[1892] = ~window[28][4];
assign temp[1893] = ~window[28][5];
assign temp[1894] = ~window[28][6];
assign temp[1895] = window[28][7];
assign temp[1896] = window[28][8];
assign temp[1920] = window[29][0];
assign temp[1921] = window[29][1];
assign temp[1922] = ~window[29][2];
assign temp[1923] = window[29][3];
assign temp[1924] = ~window[29][4];
assign temp[1925] = ~window[29][5];
assign temp[1926] = ~window[29][6];
assign temp[1927] = window[29][7];
assign temp[1928] = window[29][8];
assign temp[1952] = ~window[30][0];
assign temp[1953] = window[30][1];
assign temp[1954] = window[30][2];
assign temp[1955] = ~window[30][3];
assign temp[1956] = ~window[30][4];
assign temp[1957] = ~window[30][5];
assign temp[1958] = ~window[30][6];
assign temp[1959] = window[30][7];
assign temp[1960] = window[30][8];
assign temp[1984] = ~window[31][0];
assign temp[1985] = window[31][1];
assign temp[1986] = window[31][2];
assign temp[1987] = window[31][3];
assign temp[1988] = window[31][4];
assign temp[1989] = window[31][5];
assign temp[1990] = window[31][6];
assign temp[1991] = window[31][7];
assign temp[1992] = window[31][8];


always @(*) begin
    for (int i = 0; i < OUTPUT_CHANNELS; i++) begin
        for (int j = 0; j < INPUT_CHANNELS; j++) begin
            for (int k = 0; k < KERNEL_DIM ** 2; k++) begin
            o[i] += temp[i * OUTPUT_CHANNELS + j * INPUT_CHANNELS + k];
            end
        end
    end
end

endmodule