module classifier #(
    parameter INPUT_DIM = 784,
    parameter OUTPUT_DIM = 10
) (
    input clk,
    input reset,
    input [INPUT_DIM-1:0] inbuffer_data,
    output [$clog2(INPUT_DIM+1)+1:0] outbuffer_data,
    output reg outbuffer_we,
    output ready
);

// Enable for Icarus wavedump
// initial begin
//     $dumpfile("classifier.dmp");
//     $dumpvars();
//     // $finish();
// end

reg [$clog2(OUTPUT_DIM)-1:0] counter;

assign ready = counter == OUTPUT_DIM;

reg [INPUT_DIM-1:0] xnor_out;
wire [INPUT_DIM-1:0] xnor0;
wire [INPUT_DIM-1:0] xnor1;
wire [INPUT_DIM-1:0] xnor2;
wire [INPUT_DIM-1:0] xnor3;
wire [INPUT_DIM-1:0] xnor4;
wire [INPUT_DIM-1:0] xnor5;
wire [INPUT_DIM-1:0] xnor6;
wire [INPUT_DIM-1:0] xnor7;
wire [INPUT_DIM-1:0] xnor8;
wire [INPUT_DIM-1:0] xnor9;

// Put the other xnor outputs here as well.

// Use one popcount / activation unit for the entire layer
no_activation #(INPUT_DIM) a0 (
    .xnor_in(xnor_out),
    .logit(outbuffer_data)
);

always_ff @(posedge(clk)) begin
    if (reset) begin
        counter <= 0;
        outbuffer_we <= 1;
    end else begin
        if (counter < OUTPUT_DIM) begin
            outbuffer_we <= 1;
            counter <= counter + 1;
        end else begin
            outbuffer_we <= 0;
            counter <= counter;
        end
    end
end

always @(counter, xnor0, xnor1, xnor2, xnor3, xnor4, xnor5, xnor6, xnor7, xnor8, xnor9) begin
    case (counter)
		0 : xnor_out <= xnor0;
		1 : xnor_out <= xnor1;
		2 : xnor_out <= xnor2;
		3 : xnor_out <= xnor3;
		4 : xnor_out <= xnor4;
		5 : xnor_out <= xnor5;
		6 : xnor_out <= xnor6;
		7 : xnor_out <= xnor7;
		8 : xnor_out <= xnor8;
		9 : xnor_out <= xnor9;

        default : xnor_out <= xnor0;
    endcase
end

// Here goes the myriad of assign statements
assign xnor0[0] = 1'b1 ^~ inbuffer_data[0];
assign xnor0[1] = 1'b1 ^~ inbuffer_data[1];
assign xnor0[2] = 1'b0 ^~ inbuffer_data[2];
assign xnor0[3] = 1'b0 ^~ inbuffer_data[3];
assign xnor0[4] = 1'b0 ^~ inbuffer_data[4];
assign xnor0[5] = 1'b0 ^~ inbuffer_data[5];
assign xnor0[6] = 1'b1 ^~ inbuffer_data[6];
assign xnor0[7] = 1'b1 ^~ inbuffer_data[7];
assign xnor0[8] = 1'b1 ^~ inbuffer_data[8];
assign xnor0[9] = 1'b1 ^~ inbuffer_data[9];
assign xnor0[10] = 1'b1 ^~ inbuffer_data[10];
assign xnor0[11] = 1'b0 ^~ inbuffer_data[11];
assign xnor0[12] = 1'b1 ^~ inbuffer_data[12];
assign xnor0[13] = 1'b1 ^~ inbuffer_data[13];
assign xnor0[14] = 1'b1 ^~ inbuffer_data[14];
assign xnor0[15] = 1'b0 ^~ inbuffer_data[15];
assign xnor0[16] = 1'b1 ^~ inbuffer_data[16];
assign xnor0[17] = 1'b0 ^~ inbuffer_data[17];
assign xnor0[18] = 1'b0 ^~ inbuffer_data[18];
assign xnor0[19] = 1'b1 ^~ inbuffer_data[19];
assign xnor0[20] = 1'b1 ^~ inbuffer_data[20];
assign xnor0[21] = 1'b0 ^~ inbuffer_data[21];
assign xnor0[22] = 1'b0 ^~ inbuffer_data[22];
assign xnor0[23] = 1'b1 ^~ inbuffer_data[23];
assign xnor0[24] = 1'b1 ^~ inbuffer_data[24];
assign xnor0[25] = 1'b1 ^~ inbuffer_data[25];
assign xnor0[26] = 1'b0 ^~ inbuffer_data[26];
assign xnor0[27] = 1'b1 ^~ inbuffer_data[27];
assign xnor0[28] = 1'b0 ^~ inbuffer_data[28];
assign xnor0[29] = 1'b1 ^~ inbuffer_data[29];
assign xnor0[30] = 1'b1 ^~ inbuffer_data[30];
assign xnor0[31] = 1'b1 ^~ inbuffer_data[31];
assign xnor0[32] = 1'b1 ^~ inbuffer_data[32];
assign xnor0[33] = 1'b1 ^~ inbuffer_data[33];
assign xnor0[34] = 1'b1 ^~ inbuffer_data[34];
assign xnor0[35] = 1'b0 ^~ inbuffer_data[35];
assign xnor0[36] = 1'b0 ^~ inbuffer_data[36];
assign xnor0[37] = 1'b0 ^~ inbuffer_data[37];
assign xnor0[38] = 1'b1 ^~ inbuffer_data[38];
assign xnor0[39] = 1'b1 ^~ inbuffer_data[39];
assign xnor0[40] = 1'b0 ^~ inbuffer_data[40];
assign xnor0[41] = 1'b0 ^~ inbuffer_data[41];
assign xnor0[42] = 1'b1 ^~ inbuffer_data[42];
assign xnor0[43] = 1'b1 ^~ inbuffer_data[43];
assign xnor0[44] = 1'b0 ^~ inbuffer_data[44];
assign xnor0[45] = 1'b1 ^~ inbuffer_data[45];
assign xnor0[46] = 1'b0 ^~ inbuffer_data[46];
assign xnor0[47] = 1'b1 ^~ inbuffer_data[47];
assign xnor0[48] = 1'b0 ^~ inbuffer_data[48];
assign xnor0[49] = 1'b1 ^~ inbuffer_data[49];
assign xnor0[50] = 1'b0 ^~ inbuffer_data[50];
assign xnor0[51] = 1'b0 ^~ inbuffer_data[51];
assign xnor0[52] = 1'b0 ^~ inbuffer_data[52];
assign xnor0[53] = 1'b1 ^~ inbuffer_data[53];
assign xnor0[54] = 1'b1 ^~ inbuffer_data[54];
assign xnor0[55] = 1'b0 ^~ inbuffer_data[55];
assign xnor0[56] = 1'b0 ^~ inbuffer_data[56];
assign xnor0[57] = 1'b1 ^~ inbuffer_data[57];
assign xnor0[58] = 1'b0 ^~ inbuffer_data[58];
assign xnor0[59] = 1'b0 ^~ inbuffer_data[59];
assign xnor0[60] = 1'b1 ^~ inbuffer_data[60];
assign xnor0[61] = 1'b1 ^~ inbuffer_data[61];
assign xnor0[62] = 1'b0 ^~ inbuffer_data[62];
assign xnor0[63] = 1'b0 ^~ inbuffer_data[63];
assign xnor0[64] = 1'b0 ^~ inbuffer_data[64];
assign xnor0[65] = 1'b0 ^~ inbuffer_data[65];
assign xnor0[66] = 1'b0 ^~ inbuffer_data[66];
assign xnor0[67] = 1'b1 ^~ inbuffer_data[67];
assign xnor0[68] = 1'b1 ^~ inbuffer_data[68];
assign xnor0[69] = 1'b0 ^~ inbuffer_data[69];
assign xnor0[70] = 1'b0 ^~ inbuffer_data[70];
assign xnor0[71] = 1'b0 ^~ inbuffer_data[71];
assign xnor0[72] = 1'b1 ^~ inbuffer_data[72];
assign xnor0[73] = 1'b0 ^~ inbuffer_data[73];
assign xnor0[74] = 1'b0 ^~ inbuffer_data[74];
assign xnor0[75] = 1'b0 ^~ inbuffer_data[75];
assign xnor0[76] = 1'b1 ^~ inbuffer_data[76];
assign xnor0[77] = 1'b0 ^~ inbuffer_data[77];
assign xnor0[78] = 1'b1 ^~ inbuffer_data[78];
assign xnor0[79] = 1'b0 ^~ inbuffer_data[79];
assign xnor0[80] = 1'b0 ^~ inbuffer_data[80];
assign xnor0[81] = 1'b1 ^~ inbuffer_data[81];
assign xnor0[82] = 1'b0 ^~ inbuffer_data[82];
assign xnor0[83] = 1'b1 ^~ inbuffer_data[83];
assign xnor0[84] = 1'b0 ^~ inbuffer_data[84];
assign xnor0[85] = 1'b1 ^~ inbuffer_data[85];
assign xnor0[86] = 1'b1 ^~ inbuffer_data[86];
assign xnor0[87] = 1'b0 ^~ inbuffer_data[87];
assign xnor0[88] = 1'b1 ^~ inbuffer_data[88];
assign xnor0[89] = 1'b1 ^~ inbuffer_data[89];
assign xnor0[90] = 1'b0 ^~ inbuffer_data[90];
assign xnor0[91] = 1'b0 ^~ inbuffer_data[91];
assign xnor0[92] = 1'b0 ^~ inbuffer_data[92];
assign xnor0[93] = 1'b0 ^~ inbuffer_data[93];
assign xnor0[94] = 1'b0 ^~ inbuffer_data[94];
assign xnor0[95] = 1'b1 ^~ inbuffer_data[95];
assign xnor0[96] = 1'b0 ^~ inbuffer_data[96];
assign xnor0[97] = 1'b0 ^~ inbuffer_data[97];
assign xnor0[98] = 1'b1 ^~ inbuffer_data[98];
assign xnor0[99] = 1'b0 ^~ inbuffer_data[99];
assign xnor0[100] = 1'b0 ^~ inbuffer_data[100];
assign xnor0[101] = 1'b0 ^~ inbuffer_data[101];
assign xnor0[102] = 1'b0 ^~ inbuffer_data[102];
assign xnor0[103] = 1'b0 ^~ inbuffer_data[103];
assign xnor0[104] = 1'b0 ^~ inbuffer_data[104];
assign xnor0[105] = 1'b0 ^~ inbuffer_data[105];
assign xnor0[106] = 1'b0 ^~ inbuffer_data[106];
assign xnor0[107] = 1'b1 ^~ inbuffer_data[107];
assign xnor0[108] = 1'b0 ^~ inbuffer_data[108];
assign xnor0[109] = 1'b1 ^~ inbuffer_data[109];
assign xnor0[110] = 1'b1 ^~ inbuffer_data[110];
assign xnor0[111] = 1'b0 ^~ inbuffer_data[111];
assign xnor0[112] = 1'b0 ^~ inbuffer_data[112];
assign xnor0[113] = 1'b1 ^~ inbuffer_data[113];
assign xnor0[114] = 1'b0 ^~ inbuffer_data[114];
assign xnor0[115] = 1'b1 ^~ inbuffer_data[115];
assign xnor0[116] = 1'b1 ^~ inbuffer_data[116];
assign xnor0[117] = 1'b0 ^~ inbuffer_data[117];
assign xnor0[118] = 1'b1 ^~ inbuffer_data[118];
assign xnor0[119] = 1'b1 ^~ inbuffer_data[119];
assign xnor0[120] = 1'b0 ^~ inbuffer_data[120];
assign xnor0[121] = 1'b1 ^~ inbuffer_data[121];
assign xnor0[122] = 1'b0 ^~ inbuffer_data[122];
assign xnor0[123] = 1'b0 ^~ inbuffer_data[123];
assign xnor0[124] = 1'b0 ^~ inbuffer_data[124];
assign xnor0[125] = 1'b1 ^~ inbuffer_data[125];
assign xnor0[126] = 1'b0 ^~ inbuffer_data[126];
assign xnor0[127] = 1'b1 ^~ inbuffer_data[127];
assign xnor0[128] = 1'b1 ^~ inbuffer_data[128];
assign xnor0[129] = 1'b1 ^~ inbuffer_data[129];
assign xnor0[130] = 1'b0 ^~ inbuffer_data[130];
assign xnor0[131] = 1'b0 ^~ inbuffer_data[131];
assign xnor0[132] = 1'b0 ^~ inbuffer_data[132];
assign xnor0[133] = 1'b1 ^~ inbuffer_data[133];
assign xnor0[134] = 1'b0 ^~ inbuffer_data[134];
assign xnor0[135] = 1'b0 ^~ inbuffer_data[135];
assign xnor0[136] = 1'b0 ^~ inbuffer_data[136];
assign xnor0[137] = 1'b1 ^~ inbuffer_data[137];
assign xnor0[138] = 1'b0 ^~ inbuffer_data[138];
assign xnor0[139] = 1'b0 ^~ inbuffer_data[139];
assign xnor0[140] = 1'b1 ^~ inbuffer_data[140];
assign xnor0[141] = 1'b1 ^~ inbuffer_data[141];
assign xnor0[142] = 1'b1 ^~ inbuffer_data[142];
assign xnor0[143] = 1'b0 ^~ inbuffer_data[143];
assign xnor0[144] = 1'b0 ^~ inbuffer_data[144];
assign xnor0[145] = 1'b1 ^~ inbuffer_data[145];
assign xnor0[146] = 1'b0 ^~ inbuffer_data[146];
assign xnor0[147] = 1'b0 ^~ inbuffer_data[147];
assign xnor0[148] = 1'b1 ^~ inbuffer_data[148];
assign xnor0[149] = 1'b0 ^~ inbuffer_data[149];
assign xnor0[150] = 1'b1 ^~ inbuffer_data[150];
assign xnor0[151] = 1'b1 ^~ inbuffer_data[151];
assign xnor0[152] = 1'b1 ^~ inbuffer_data[152];
assign xnor0[153] = 1'b1 ^~ inbuffer_data[153];
assign xnor0[154] = 1'b1 ^~ inbuffer_data[154];
assign xnor0[155] = 1'b1 ^~ inbuffer_data[155];
assign xnor0[156] = 1'b1 ^~ inbuffer_data[156];
assign xnor0[157] = 1'b1 ^~ inbuffer_data[157];
assign xnor0[158] = 1'b1 ^~ inbuffer_data[158];
assign xnor0[159] = 1'b0 ^~ inbuffer_data[159];
assign xnor0[160] = 1'b0 ^~ inbuffer_data[160];
assign xnor0[161] = 1'b0 ^~ inbuffer_data[161];
assign xnor0[162] = 1'b1 ^~ inbuffer_data[162];
assign xnor0[163] = 1'b0 ^~ inbuffer_data[163];
assign xnor0[164] = 1'b0 ^~ inbuffer_data[164];
assign xnor0[165] = 1'b0 ^~ inbuffer_data[165];
assign xnor0[166] = 1'b1 ^~ inbuffer_data[166];
assign xnor0[167] = 1'b0 ^~ inbuffer_data[167];
assign xnor0[168] = 1'b0 ^~ inbuffer_data[168];
assign xnor0[169] = 1'b1 ^~ inbuffer_data[169];
assign xnor0[170] = 1'b1 ^~ inbuffer_data[170];
assign xnor0[171] = 1'b1 ^~ inbuffer_data[171];
assign xnor0[172] = 1'b0 ^~ inbuffer_data[172];
assign xnor0[173] = 1'b0 ^~ inbuffer_data[173];
assign xnor0[174] = 1'b0 ^~ inbuffer_data[174];
assign xnor0[175] = 1'b0 ^~ inbuffer_data[175];
assign xnor0[176] = 1'b0 ^~ inbuffer_data[176];
assign xnor0[177] = 1'b0 ^~ inbuffer_data[177];
assign xnor0[178] = 1'b0 ^~ inbuffer_data[178];
assign xnor0[179] = 1'b0 ^~ inbuffer_data[179];
assign xnor0[180] = 1'b1 ^~ inbuffer_data[180];
assign xnor0[181] = 1'b0 ^~ inbuffer_data[181];
assign xnor0[182] = 1'b0 ^~ inbuffer_data[182];
assign xnor0[183] = 1'b1 ^~ inbuffer_data[183];
assign xnor0[184] = 1'b1 ^~ inbuffer_data[184];
assign xnor0[185] = 1'b1 ^~ inbuffer_data[185];
assign xnor0[186] = 1'b1 ^~ inbuffer_data[186];
assign xnor0[187] = 1'b1 ^~ inbuffer_data[187];
assign xnor0[188] = 1'b1 ^~ inbuffer_data[188];
assign xnor0[189] = 1'b1 ^~ inbuffer_data[189];
assign xnor0[190] = 1'b0 ^~ inbuffer_data[190];
assign xnor0[191] = 1'b0 ^~ inbuffer_data[191];
assign xnor0[192] = 1'b0 ^~ inbuffer_data[192];
assign xnor0[193] = 1'b0 ^~ inbuffer_data[193];
assign xnor0[194] = 1'b1 ^~ inbuffer_data[194];
assign xnor0[195] = 1'b0 ^~ inbuffer_data[195];
assign xnor0[196] = 1'b0 ^~ inbuffer_data[196];
assign xnor0[197] = 1'b1 ^~ inbuffer_data[197];
assign xnor0[198] = 1'b1 ^~ inbuffer_data[198];
assign xnor0[199] = 1'b1 ^~ inbuffer_data[199];
assign xnor0[200] = 1'b0 ^~ inbuffer_data[200];
assign xnor0[201] = 1'b1 ^~ inbuffer_data[201];
assign xnor0[202] = 1'b1 ^~ inbuffer_data[202];
assign xnor0[203] = 1'b1 ^~ inbuffer_data[203];
assign xnor0[204] = 1'b0 ^~ inbuffer_data[204];
assign xnor0[205] = 1'b0 ^~ inbuffer_data[205];
assign xnor0[206] = 1'b0 ^~ inbuffer_data[206];
assign xnor0[207] = 1'b1 ^~ inbuffer_data[207];
assign xnor0[208] = 1'b1 ^~ inbuffer_data[208];
assign xnor0[209] = 1'b0 ^~ inbuffer_data[209];
assign xnor0[210] = 1'b0 ^~ inbuffer_data[210];
assign xnor0[211] = 1'b1 ^~ inbuffer_data[211];
assign xnor0[212] = 1'b0 ^~ inbuffer_data[212];
assign xnor0[213] = 1'b1 ^~ inbuffer_data[213];
assign xnor0[214] = 1'b1 ^~ inbuffer_data[214];
assign xnor0[215] = 1'b1 ^~ inbuffer_data[215];
assign xnor0[216] = 1'b0 ^~ inbuffer_data[216];
assign xnor0[217] = 1'b1 ^~ inbuffer_data[217];
assign xnor0[218] = 1'b1 ^~ inbuffer_data[218];
assign xnor0[219] = 1'b1 ^~ inbuffer_data[219];
assign xnor0[220] = 1'b0 ^~ inbuffer_data[220];
assign xnor0[221] = 1'b0 ^~ inbuffer_data[221];
assign xnor0[222] = 1'b0 ^~ inbuffer_data[222];
assign xnor0[223] = 1'b0 ^~ inbuffer_data[223];
assign xnor0[224] = 1'b0 ^~ inbuffer_data[224];
assign xnor0[225] = 1'b1 ^~ inbuffer_data[225];
assign xnor0[226] = 1'b0 ^~ inbuffer_data[226];
assign xnor0[227] = 1'b0 ^~ inbuffer_data[227];
assign xnor0[228] = 1'b0 ^~ inbuffer_data[228];
assign xnor0[229] = 1'b1 ^~ inbuffer_data[229];
assign xnor0[230] = 1'b0 ^~ inbuffer_data[230];
assign xnor0[231] = 1'b0 ^~ inbuffer_data[231];
assign xnor0[232] = 1'b1 ^~ inbuffer_data[232];
assign xnor0[233] = 1'b1 ^~ inbuffer_data[233];
assign xnor0[234] = 1'b1 ^~ inbuffer_data[234];
assign xnor0[235] = 1'b1 ^~ inbuffer_data[235];
assign xnor0[236] = 1'b1 ^~ inbuffer_data[236];
assign xnor0[237] = 1'b1 ^~ inbuffer_data[237];
assign xnor0[238] = 1'b1 ^~ inbuffer_data[238];
assign xnor0[239] = 1'b1 ^~ inbuffer_data[239];
assign xnor0[240] = 1'b1 ^~ inbuffer_data[240];
assign xnor0[241] = 1'b1 ^~ inbuffer_data[241];
assign xnor0[242] = 1'b1 ^~ inbuffer_data[242];
assign xnor0[243] = 1'b1 ^~ inbuffer_data[243];
assign xnor0[244] = 1'b0 ^~ inbuffer_data[244];
assign xnor0[245] = 1'b1 ^~ inbuffer_data[245];
assign xnor0[246] = 1'b0 ^~ inbuffer_data[246];
assign xnor0[247] = 1'b1 ^~ inbuffer_data[247];
assign xnor0[248] = 1'b0 ^~ inbuffer_data[248];
assign xnor0[249] = 1'b0 ^~ inbuffer_data[249];
assign xnor0[250] = 1'b0 ^~ inbuffer_data[250];
assign xnor0[251] = 1'b1 ^~ inbuffer_data[251];
assign xnor0[252] = 1'b1 ^~ inbuffer_data[252];
assign xnor0[253] = 1'b0 ^~ inbuffer_data[253];
assign xnor0[254] = 1'b1 ^~ inbuffer_data[254];
assign xnor0[255] = 1'b0 ^~ inbuffer_data[255];
assign xnor0[256] = 1'b0 ^~ inbuffer_data[256];
assign xnor0[257] = 1'b0 ^~ inbuffer_data[257];
assign xnor0[258] = 1'b0 ^~ inbuffer_data[258];
assign xnor0[259] = 1'b1 ^~ inbuffer_data[259];
assign xnor0[260] = 1'b0 ^~ inbuffer_data[260];
assign xnor0[261] = 1'b0 ^~ inbuffer_data[261];
assign xnor0[262] = 1'b1 ^~ inbuffer_data[262];
assign xnor0[263] = 1'b1 ^~ inbuffer_data[263];
assign xnor0[264] = 1'b1 ^~ inbuffer_data[264];
assign xnor0[265] = 1'b1 ^~ inbuffer_data[265];
assign xnor0[266] = 1'b1 ^~ inbuffer_data[266];
assign xnor0[267] = 1'b0 ^~ inbuffer_data[267];
assign xnor0[268] = 1'b1 ^~ inbuffer_data[268];
assign xnor0[269] = 1'b1 ^~ inbuffer_data[269];
assign xnor0[270] = 1'b1 ^~ inbuffer_data[270];
assign xnor0[271] = 1'b1 ^~ inbuffer_data[271];
assign xnor0[272] = 1'b0 ^~ inbuffer_data[272];
assign xnor0[273] = 1'b0 ^~ inbuffer_data[273];
assign xnor0[274] = 1'b1 ^~ inbuffer_data[274];
assign xnor0[275] = 1'b1 ^~ inbuffer_data[275];
assign xnor0[276] = 1'b0 ^~ inbuffer_data[276];
assign xnor0[277] = 1'b0 ^~ inbuffer_data[277];
assign xnor0[278] = 1'b0 ^~ inbuffer_data[278];
assign xnor0[279] = 1'b1 ^~ inbuffer_data[279];
assign xnor0[280] = 1'b0 ^~ inbuffer_data[280];
assign xnor0[281] = 1'b1 ^~ inbuffer_data[281];
assign xnor0[282] = 1'b1 ^~ inbuffer_data[282];
assign xnor0[283] = 1'b1 ^~ inbuffer_data[283];
assign xnor0[284] = 1'b1 ^~ inbuffer_data[284];
assign xnor0[285] = 1'b1 ^~ inbuffer_data[285];
assign xnor0[286] = 1'b0 ^~ inbuffer_data[286];
assign xnor0[287] = 1'b0 ^~ inbuffer_data[287];
assign xnor0[288] = 1'b0 ^~ inbuffer_data[288];
assign xnor0[289] = 1'b0 ^~ inbuffer_data[289];
assign xnor0[290] = 1'b0 ^~ inbuffer_data[290];
assign xnor0[291] = 1'b1 ^~ inbuffer_data[291];
assign xnor0[292] = 1'b1 ^~ inbuffer_data[292];
assign xnor0[293] = 1'b0 ^~ inbuffer_data[293];
assign xnor0[294] = 1'b1 ^~ inbuffer_data[294];
assign xnor0[295] = 1'b0 ^~ inbuffer_data[295];
assign xnor0[296] = 1'b0 ^~ inbuffer_data[296];
assign xnor0[297] = 1'b1 ^~ inbuffer_data[297];
assign xnor0[298] = 1'b1 ^~ inbuffer_data[298];
assign xnor0[299] = 1'b1 ^~ inbuffer_data[299];
assign xnor0[300] = 1'b1 ^~ inbuffer_data[300];
assign xnor0[301] = 1'b1 ^~ inbuffer_data[301];
assign xnor0[302] = 1'b1 ^~ inbuffer_data[302];
assign xnor0[303] = 1'b1 ^~ inbuffer_data[303];
assign xnor0[304] = 1'b0 ^~ inbuffer_data[304];
assign xnor0[305] = 1'b0 ^~ inbuffer_data[305];
assign xnor0[306] = 1'b0 ^~ inbuffer_data[306];
assign xnor0[307] = 1'b0 ^~ inbuffer_data[307];
assign xnor0[308] = 1'b1 ^~ inbuffer_data[308];
assign xnor0[309] = 1'b0 ^~ inbuffer_data[309];
assign xnor0[310] = 1'b0 ^~ inbuffer_data[310];
assign xnor0[311] = 1'b0 ^~ inbuffer_data[311];
assign xnor0[312] = 1'b0 ^~ inbuffer_data[312];
assign xnor0[313] = 1'b0 ^~ inbuffer_data[313];
assign xnor0[314] = 1'b1 ^~ inbuffer_data[314];
assign xnor0[315] = 1'b1 ^~ inbuffer_data[315];
assign xnor0[316] = 1'b1 ^~ inbuffer_data[316];
assign xnor0[317] = 1'b0 ^~ inbuffer_data[317];
assign xnor0[318] = 1'b0 ^~ inbuffer_data[318];
assign xnor0[319] = 1'b0 ^~ inbuffer_data[319];
assign xnor0[320] = 1'b0 ^~ inbuffer_data[320];
assign xnor0[321] = 1'b0 ^~ inbuffer_data[321];
assign xnor0[322] = 1'b0 ^~ inbuffer_data[322];
assign xnor0[323] = 1'b0 ^~ inbuffer_data[323];
assign xnor0[324] = 1'b0 ^~ inbuffer_data[324];
assign xnor0[325] = 1'b0 ^~ inbuffer_data[325];
assign xnor0[326] = 1'b0 ^~ inbuffer_data[326];
assign xnor0[327] = 1'b1 ^~ inbuffer_data[327];
assign xnor0[328] = 1'b1 ^~ inbuffer_data[328];
assign xnor0[329] = 1'b1 ^~ inbuffer_data[329];
assign xnor0[330] = 1'b1 ^~ inbuffer_data[330];
assign xnor0[331] = 1'b1 ^~ inbuffer_data[331];
assign xnor0[332] = 1'b1 ^~ inbuffer_data[332];
assign xnor0[333] = 1'b0 ^~ inbuffer_data[333];
assign xnor0[334] = 1'b0 ^~ inbuffer_data[334];
assign xnor0[335] = 1'b1 ^~ inbuffer_data[335];
assign xnor0[336] = 1'b0 ^~ inbuffer_data[336];
assign xnor0[337] = 1'b0 ^~ inbuffer_data[337];
assign xnor0[338] = 1'b0 ^~ inbuffer_data[338];
assign xnor0[339] = 1'b0 ^~ inbuffer_data[339];
assign xnor0[340] = 1'b0 ^~ inbuffer_data[340];
assign xnor0[341] = 1'b1 ^~ inbuffer_data[341];
assign xnor0[342] = 1'b1 ^~ inbuffer_data[342];
assign xnor0[343] = 1'b1 ^~ inbuffer_data[343];
assign xnor0[344] = 1'b0 ^~ inbuffer_data[344];
assign xnor0[345] = 1'b1 ^~ inbuffer_data[345];
assign xnor0[346] = 1'b1 ^~ inbuffer_data[346];
assign xnor0[347] = 1'b0 ^~ inbuffer_data[347];
assign xnor0[348] = 1'b1 ^~ inbuffer_data[348];
assign xnor0[349] = 1'b0 ^~ inbuffer_data[349];
assign xnor0[350] = 1'b0 ^~ inbuffer_data[350];
assign xnor0[351] = 1'b0 ^~ inbuffer_data[351];
assign xnor0[352] = 1'b0 ^~ inbuffer_data[352];
assign xnor0[353] = 1'b0 ^~ inbuffer_data[353];
assign xnor0[354] = 1'b0 ^~ inbuffer_data[354];
assign xnor0[355] = 1'b0 ^~ inbuffer_data[355];
assign xnor0[356] = 1'b0 ^~ inbuffer_data[356];
assign xnor0[357] = 1'b1 ^~ inbuffer_data[357];
assign xnor0[358] = 1'b1 ^~ inbuffer_data[358];
assign xnor0[359] = 1'b1 ^~ inbuffer_data[359];
assign xnor0[360] = 1'b1 ^~ inbuffer_data[360];
assign xnor0[361] = 1'b1 ^~ inbuffer_data[361];
assign xnor0[362] = 1'b0 ^~ inbuffer_data[362];
assign xnor0[363] = 1'b1 ^~ inbuffer_data[363];
assign xnor0[364] = 1'b0 ^~ inbuffer_data[364];
assign xnor0[365] = 1'b1 ^~ inbuffer_data[365];
assign xnor0[366] = 1'b1 ^~ inbuffer_data[366];
assign xnor0[367] = 1'b1 ^~ inbuffer_data[367];
assign xnor0[368] = 1'b0 ^~ inbuffer_data[368];
assign xnor0[369] = 1'b1 ^~ inbuffer_data[369];
assign xnor0[370] = 1'b1 ^~ inbuffer_data[370];
assign xnor0[371] = 1'b1 ^~ inbuffer_data[371];
assign xnor0[372] = 1'b1 ^~ inbuffer_data[372];
assign xnor0[373] = 1'b1 ^~ inbuffer_data[373];
assign xnor0[374] = 1'b1 ^~ inbuffer_data[374];
assign xnor0[375] = 1'b1 ^~ inbuffer_data[375];
assign xnor0[376] = 1'b0 ^~ inbuffer_data[376];
assign xnor0[377] = 1'b0 ^~ inbuffer_data[377];
assign xnor0[378] = 1'b0 ^~ inbuffer_data[378];
assign xnor0[379] = 1'b0 ^~ inbuffer_data[379];
assign xnor0[380] = 1'b0 ^~ inbuffer_data[380];
assign xnor0[381] = 1'b0 ^~ inbuffer_data[381];
assign xnor0[382] = 1'b0 ^~ inbuffer_data[382];
assign xnor0[383] = 1'b0 ^~ inbuffer_data[383];
assign xnor0[384] = 1'b0 ^~ inbuffer_data[384];
assign xnor0[385] = 1'b1 ^~ inbuffer_data[385];
assign xnor0[386] = 1'b1 ^~ inbuffer_data[386];
assign xnor0[387] = 1'b1 ^~ inbuffer_data[387];
assign xnor0[388] = 1'b1 ^~ inbuffer_data[388];
assign xnor0[389] = 1'b0 ^~ inbuffer_data[389];
assign xnor0[390] = 1'b1 ^~ inbuffer_data[390];
assign xnor0[391] = 1'b1 ^~ inbuffer_data[391];
assign xnor0[392] = 1'b1 ^~ inbuffer_data[392];
assign xnor0[393] = 1'b0 ^~ inbuffer_data[393];
assign xnor0[394] = 1'b0 ^~ inbuffer_data[394];
assign xnor0[395] = 1'b0 ^~ inbuffer_data[395];
assign xnor0[396] = 1'b1 ^~ inbuffer_data[396];
assign xnor0[397] = 1'b1 ^~ inbuffer_data[397];
assign xnor0[398] = 1'b1 ^~ inbuffer_data[398];
assign xnor0[399] = 1'b1 ^~ inbuffer_data[399];
assign xnor0[400] = 1'b1 ^~ inbuffer_data[400];
assign xnor0[401] = 1'b1 ^~ inbuffer_data[401];
assign xnor0[402] = 1'b0 ^~ inbuffer_data[402];
assign xnor0[403] = 1'b1 ^~ inbuffer_data[403];
assign xnor0[404] = 1'b0 ^~ inbuffer_data[404];
assign xnor0[405] = 1'b0 ^~ inbuffer_data[405];
assign xnor0[406] = 1'b0 ^~ inbuffer_data[406];
assign xnor0[407] = 1'b0 ^~ inbuffer_data[407];
assign xnor0[408] = 1'b0 ^~ inbuffer_data[408];
assign xnor0[409] = 1'b0 ^~ inbuffer_data[409];
assign xnor0[410] = 1'b0 ^~ inbuffer_data[410];
assign xnor0[411] = 1'b0 ^~ inbuffer_data[411];
assign xnor0[412] = 1'b1 ^~ inbuffer_data[412];
assign xnor0[413] = 1'b1 ^~ inbuffer_data[413];
assign xnor0[414] = 1'b1 ^~ inbuffer_data[414];
assign xnor0[415] = 1'b1 ^~ inbuffer_data[415];
assign xnor0[416] = 1'b1 ^~ inbuffer_data[416];
assign xnor0[417] = 1'b0 ^~ inbuffer_data[417];
assign xnor0[418] = 1'b1 ^~ inbuffer_data[418];
assign xnor0[419] = 1'b0 ^~ inbuffer_data[419];
assign xnor0[420] = 1'b0 ^~ inbuffer_data[420];
assign xnor0[421] = 1'b1 ^~ inbuffer_data[421];
assign xnor0[422] = 1'b0 ^~ inbuffer_data[422];
assign xnor0[423] = 1'b1 ^~ inbuffer_data[423];
assign xnor0[424] = 1'b1 ^~ inbuffer_data[424];
assign xnor0[425] = 1'b1 ^~ inbuffer_data[425];
assign xnor0[426] = 1'b1 ^~ inbuffer_data[426];
assign xnor0[427] = 1'b1 ^~ inbuffer_data[427];
assign xnor0[428] = 1'b1 ^~ inbuffer_data[428];
assign xnor0[429] = 1'b1 ^~ inbuffer_data[429];
assign xnor0[430] = 1'b1 ^~ inbuffer_data[430];
assign xnor0[431] = 1'b1 ^~ inbuffer_data[431];
assign xnor0[432] = 1'b0 ^~ inbuffer_data[432];
assign xnor0[433] = 1'b0 ^~ inbuffer_data[433];
assign xnor0[434] = 1'b0 ^~ inbuffer_data[434];
assign xnor0[435] = 1'b0 ^~ inbuffer_data[435];
assign xnor0[436] = 1'b0 ^~ inbuffer_data[436];
assign xnor0[437] = 1'b0 ^~ inbuffer_data[437];
assign xnor0[438] = 1'b0 ^~ inbuffer_data[438];
assign xnor0[439] = 1'b1 ^~ inbuffer_data[439];
assign xnor0[440] = 1'b1 ^~ inbuffer_data[440];
assign xnor0[441] = 1'b1 ^~ inbuffer_data[441];
assign xnor0[442] = 1'b1 ^~ inbuffer_data[442];
assign xnor0[443] = 1'b1 ^~ inbuffer_data[443];
assign xnor0[444] = 1'b1 ^~ inbuffer_data[444];
assign xnor0[445] = 1'b1 ^~ inbuffer_data[445];
assign xnor0[446] = 1'b0 ^~ inbuffer_data[446];
assign xnor0[447] = 1'b1 ^~ inbuffer_data[447];
assign xnor0[448] = 1'b1 ^~ inbuffer_data[448];
assign xnor0[449] = 1'b0 ^~ inbuffer_data[449];
assign xnor0[450] = 1'b0 ^~ inbuffer_data[450];
assign xnor0[451] = 1'b0 ^~ inbuffer_data[451];
assign xnor0[452] = 1'b0 ^~ inbuffer_data[452];
assign xnor0[453] = 1'b1 ^~ inbuffer_data[453];
assign xnor0[454] = 1'b1 ^~ inbuffer_data[454];
assign xnor0[455] = 1'b1 ^~ inbuffer_data[455];
assign xnor0[456] = 1'b1 ^~ inbuffer_data[456];
assign xnor0[457] = 1'b1 ^~ inbuffer_data[457];
assign xnor0[458] = 1'b1 ^~ inbuffer_data[458];
assign xnor0[459] = 1'b0 ^~ inbuffer_data[459];
assign xnor0[460] = 1'b0 ^~ inbuffer_data[460];
assign xnor0[461] = 1'b0 ^~ inbuffer_data[461];
assign xnor0[462] = 1'b0 ^~ inbuffer_data[462];
assign xnor0[463] = 1'b0 ^~ inbuffer_data[463];
assign xnor0[464] = 1'b0 ^~ inbuffer_data[464];
assign xnor0[465] = 1'b0 ^~ inbuffer_data[465];
assign xnor0[466] = 1'b1 ^~ inbuffer_data[466];
assign xnor0[467] = 1'b0 ^~ inbuffer_data[467];
assign xnor0[468] = 1'b1 ^~ inbuffer_data[468];
assign xnor0[469] = 1'b1 ^~ inbuffer_data[469];
assign xnor0[470] = 1'b1 ^~ inbuffer_data[470];
assign xnor0[471] = 1'b1 ^~ inbuffer_data[471];
assign xnor0[472] = 1'b1 ^~ inbuffer_data[472];
assign xnor0[473] = 1'b0 ^~ inbuffer_data[473];
assign xnor0[474] = 1'b0 ^~ inbuffer_data[474];
assign xnor0[475] = 1'b1 ^~ inbuffer_data[475];
assign xnor0[476] = 1'b1 ^~ inbuffer_data[476];
assign xnor0[477] = 1'b1 ^~ inbuffer_data[477];
assign xnor0[478] = 1'b0 ^~ inbuffer_data[478];
assign xnor0[479] = 1'b0 ^~ inbuffer_data[479];
assign xnor0[480] = 1'b0 ^~ inbuffer_data[480];
assign xnor0[481] = 1'b1 ^~ inbuffer_data[481];
assign xnor0[482] = 1'b1 ^~ inbuffer_data[482];
assign xnor0[483] = 1'b1 ^~ inbuffer_data[483];
assign xnor0[484] = 1'b1 ^~ inbuffer_data[484];
assign xnor0[485] = 1'b1 ^~ inbuffer_data[485];
assign xnor0[486] = 1'b1 ^~ inbuffer_data[486];
assign xnor0[487] = 1'b0 ^~ inbuffer_data[487];
assign xnor0[488] = 1'b0 ^~ inbuffer_data[488];
assign xnor0[489] = 1'b0 ^~ inbuffer_data[489];
assign xnor0[490] = 1'b0 ^~ inbuffer_data[490];
assign xnor0[491] = 1'b0 ^~ inbuffer_data[491];
assign xnor0[492] = 1'b0 ^~ inbuffer_data[492];
assign xnor0[493] = 1'b1 ^~ inbuffer_data[493];
assign xnor0[494] = 1'b1 ^~ inbuffer_data[494];
assign xnor0[495] = 1'b0 ^~ inbuffer_data[495];
assign xnor0[496] = 1'b0 ^~ inbuffer_data[496];
assign xnor0[497] = 1'b0 ^~ inbuffer_data[497];
assign xnor0[498] = 1'b1 ^~ inbuffer_data[498];
assign xnor0[499] = 1'b1 ^~ inbuffer_data[499];
assign xnor0[500] = 1'b1 ^~ inbuffer_data[500];
assign xnor0[501] = 1'b1 ^~ inbuffer_data[501];
assign xnor0[502] = 1'b1 ^~ inbuffer_data[502];
assign xnor0[503] = 1'b0 ^~ inbuffer_data[503];
assign xnor0[504] = 1'b0 ^~ inbuffer_data[504];
assign xnor0[505] = 1'b0 ^~ inbuffer_data[505];
assign xnor0[506] = 1'b0 ^~ inbuffer_data[506];
assign xnor0[507] = 1'b1 ^~ inbuffer_data[507];
assign xnor0[508] = 1'b0 ^~ inbuffer_data[508];
assign xnor0[509] = 1'b1 ^~ inbuffer_data[509];
assign xnor0[510] = 1'b1 ^~ inbuffer_data[510];
assign xnor0[511] = 1'b1 ^~ inbuffer_data[511];
assign xnor0[512] = 1'b1 ^~ inbuffer_data[512];
assign xnor0[513] = 1'b1 ^~ inbuffer_data[513];
assign xnor0[514] = 1'b1 ^~ inbuffer_data[514];
assign xnor0[515] = 1'b1 ^~ inbuffer_data[515];
assign xnor0[516] = 1'b0 ^~ inbuffer_data[516];
assign xnor0[517] = 1'b0 ^~ inbuffer_data[517];
assign xnor0[518] = 1'b0 ^~ inbuffer_data[518];
assign xnor0[519] = 1'b0 ^~ inbuffer_data[519];
assign xnor0[520] = 1'b1 ^~ inbuffer_data[520];
assign xnor0[521] = 1'b1 ^~ inbuffer_data[521];
assign xnor0[522] = 1'b0 ^~ inbuffer_data[522];
assign xnor0[523] = 1'b1 ^~ inbuffer_data[523];
assign xnor0[524] = 1'b0 ^~ inbuffer_data[524];
assign xnor0[525] = 1'b0 ^~ inbuffer_data[525];
assign xnor0[526] = 1'b1 ^~ inbuffer_data[526];
assign xnor0[527] = 1'b0 ^~ inbuffer_data[527];
assign xnor0[528] = 1'b0 ^~ inbuffer_data[528];
assign xnor0[529] = 1'b1 ^~ inbuffer_data[529];
assign xnor0[530] = 1'b1 ^~ inbuffer_data[530];
assign xnor0[531] = 1'b0 ^~ inbuffer_data[531];
assign xnor0[532] = 1'b0 ^~ inbuffer_data[532];
assign xnor0[533] = 1'b0 ^~ inbuffer_data[533];
assign xnor0[534] = 1'b0 ^~ inbuffer_data[534];
assign xnor0[535] = 1'b0 ^~ inbuffer_data[535];
assign xnor0[536] = 1'b0 ^~ inbuffer_data[536];
assign xnor0[537] = 1'b1 ^~ inbuffer_data[537];
assign xnor0[538] = 1'b1 ^~ inbuffer_data[538];
assign xnor0[539] = 1'b1 ^~ inbuffer_data[539];
assign xnor0[540] = 1'b1 ^~ inbuffer_data[540];
assign xnor0[541] = 1'b1 ^~ inbuffer_data[541];
assign xnor0[542] = 1'b1 ^~ inbuffer_data[542];
assign xnor0[543] = 1'b1 ^~ inbuffer_data[543];
assign xnor0[544] = 1'b0 ^~ inbuffer_data[544];
assign xnor0[545] = 1'b0 ^~ inbuffer_data[545];
assign xnor0[546] = 1'b0 ^~ inbuffer_data[546];
assign xnor0[547] = 1'b0 ^~ inbuffer_data[547];
assign xnor0[548] = 1'b1 ^~ inbuffer_data[548];
assign xnor0[549] = 1'b1 ^~ inbuffer_data[549];
assign xnor0[550] = 1'b1 ^~ inbuffer_data[550];
assign xnor0[551] = 1'b0 ^~ inbuffer_data[551];
assign xnor0[552] = 1'b1 ^~ inbuffer_data[552];
assign xnor0[553] = 1'b0 ^~ inbuffer_data[553];
assign xnor0[554] = 1'b1 ^~ inbuffer_data[554];
assign xnor0[555] = 1'b1 ^~ inbuffer_data[555];
assign xnor0[556] = 1'b0 ^~ inbuffer_data[556];
assign xnor0[557] = 1'b1 ^~ inbuffer_data[557];
assign xnor0[558] = 1'b0 ^~ inbuffer_data[558];
assign xnor0[559] = 1'b0 ^~ inbuffer_data[559];
assign xnor0[560] = 1'b0 ^~ inbuffer_data[560];
assign xnor0[561] = 1'b1 ^~ inbuffer_data[561];
assign xnor0[562] = 1'b0 ^~ inbuffer_data[562];
assign xnor0[563] = 1'b0 ^~ inbuffer_data[563];
assign xnor0[564] = 1'b0 ^~ inbuffer_data[564];
assign xnor0[565] = 1'b1 ^~ inbuffer_data[565];
assign xnor0[566] = 1'b0 ^~ inbuffer_data[566];
assign xnor0[567] = 1'b1 ^~ inbuffer_data[567];
assign xnor0[568] = 1'b1 ^~ inbuffer_data[568];
assign xnor0[569] = 1'b1 ^~ inbuffer_data[569];
assign xnor0[570] = 1'b1 ^~ inbuffer_data[570];
assign xnor0[571] = 1'b1 ^~ inbuffer_data[571];
assign xnor0[572] = 1'b1 ^~ inbuffer_data[572];
assign xnor0[573] = 1'b1 ^~ inbuffer_data[573];
assign xnor0[574] = 1'b0 ^~ inbuffer_data[574];
assign xnor0[575] = 1'b1 ^~ inbuffer_data[575];
assign xnor0[576] = 1'b0 ^~ inbuffer_data[576];
assign xnor0[577] = 1'b0 ^~ inbuffer_data[577];
assign xnor0[578] = 1'b1 ^~ inbuffer_data[578];
assign xnor0[579] = 1'b0 ^~ inbuffer_data[579];
assign xnor0[580] = 1'b0 ^~ inbuffer_data[580];
assign xnor0[581] = 1'b1 ^~ inbuffer_data[581];
assign xnor0[582] = 1'b0 ^~ inbuffer_data[582];
assign xnor0[583] = 1'b0 ^~ inbuffer_data[583];
assign xnor0[584] = 1'b0 ^~ inbuffer_data[584];
assign xnor0[585] = 1'b0 ^~ inbuffer_data[585];
assign xnor0[586] = 1'b0 ^~ inbuffer_data[586];
assign xnor0[587] = 1'b0 ^~ inbuffer_data[587];
assign xnor0[588] = 1'b0 ^~ inbuffer_data[588];
assign xnor0[589] = 1'b1 ^~ inbuffer_data[589];
assign xnor0[590] = 1'b1 ^~ inbuffer_data[590];
assign xnor0[591] = 1'b1 ^~ inbuffer_data[591];
assign xnor0[592] = 1'b0 ^~ inbuffer_data[592];
assign xnor0[593] = 1'b1 ^~ inbuffer_data[593];
assign xnor0[594] = 1'b1 ^~ inbuffer_data[594];
assign xnor0[595] = 1'b1 ^~ inbuffer_data[595];
assign xnor0[596] = 1'b0 ^~ inbuffer_data[596];
assign xnor0[597] = 1'b1 ^~ inbuffer_data[597];
assign xnor0[598] = 1'b1 ^~ inbuffer_data[598];
assign xnor0[599] = 1'b1 ^~ inbuffer_data[599];
assign xnor0[600] = 1'b1 ^~ inbuffer_data[600];
assign xnor0[601] = 1'b1 ^~ inbuffer_data[601];
assign xnor0[602] = 1'b0 ^~ inbuffer_data[602];
assign xnor0[603] = 1'b1 ^~ inbuffer_data[603];
assign xnor0[604] = 1'b0 ^~ inbuffer_data[604];
assign xnor0[605] = 1'b0 ^~ inbuffer_data[605];
assign xnor0[606] = 1'b0 ^~ inbuffer_data[606];
assign xnor0[607] = 1'b0 ^~ inbuffer_data[607];
assign xnor0[608] = 1'b0 ^~ inbuffer_data[608];
assign xnor0[609] = 1'b0 ^~ inbuffer_data[609];
assign xnor0[610] = 1'b0 ^~ inbuffer_data[610];
assign xnor0[611] = 1'b0 ^~ inbuffer_data[611];
assign xnor0[612] = 1'b0 ^~ inbuffer_data[612];
assign xnor0[613] = 1'b1 ^~ inbuffer_data[613];
assign xnor0[614] = 1'b1 ^~ inbuffer_data[614];
assign xnor0[615] = 1'b1 ^~ inbuffer_data[615];
assign xnor0[616] = 1'b0 ^~ inbuffer_data[616];
assign xnor0[617] = 1'b1 ^~ inbuffer_data[617];
assign xnor0[618] = 1'b1 ^~ inbuffer_data[618];
assign xnor0[619] = 1'b1 ^~ inbuffer_data[619];
assign xnor0[620] = 1'b0 ^~ inbuffer_data[620];
assign xnor0[621] = 1'b0 ^~ inbuffer_data[621];
assign xnor0[622] = 1'b1 ^~ inbuffer_data[622];
assign xnor0[623] = 1'b1 ^~ inbuffer_data[623];
assign xnor0[624] = 1'b1 ^~ inbuffer_data[624];
assign xnor0[625] = 1'b1 ^~ inbuffer_data[625];
assign xnor0[626] = 1'b1 ^~ inbuffer_data[626];
assign xnor0[627] = 1'b1 ^~ inbuffer_data[627];
assign xnor0[628] = 1'b1 ^~ inbuffer_data[628];
assign xnor0[629] = 1'b1 ^~ inbuffer_data[629];
assign xnor0[630] = 1'b1 ^~ inbuffer_data[630];
assign xnor0[631] = 1'b0 ^~ inbuffer_data[631];
assign xnor0[632] = 1'b1 ^~ inbuffer_data[632];
assign xnor0[633] = 1'b0 ^~ inbuffer_data[633];
assign xnor0[634] = 1'b1 ^~ inbuffer_data[634];
assign xnor0[635] = 1'b1 ^~ inbuffer_data[635];
assign xnor0[636] = 1'b1 ^~ inbuffer_data[636];
assign xnor0[637] = 1'b0 ^~ inbuffer_data[637];
assign xnor0[638] = 1'b1 ^~ inbuffer_data[638];
assign xnor0[639] = 1'b0 ^~ inbuffer_data[639];
assign xnor0[640] = 1'b1 ^~ inbuffer_data[640];
assign xnor0[641] = 1'b0 ^~ inbuffer_data[641];
assign xnor0[642] = 1'b1 ^~ inbuffer_data[642];
assign xnor0[643] = 1'b1 ^~ inbuffer_data[643];
assign xnor0[644] = 1'b0 ^~ inbuffer_data[644];
assign xnor0[645] = 1'b0 ^~ inbuffer_data[645];
assign xnor0[646] = 1'b1 ^~ inbuffer_data[646];
assign xnor0[647] = 1'b0 ^~ inbuffer_data[647];
assign xnor0[648] = 1'b0 ^~ inbuffer_data[648];
assign xnor0[649] = 1'b0 ^~ inbuffer_data[649];
assign xnor0[650] = 1'b0 ^~ inbuffer_data[650];
assign xnor0[651] = 1'b1 ^~ inbuffer_data[651];
assign xnor0[652] = 1'b1 ^~ inbuffer_data[652];
assign xnor0[653] = 1'b1 ^~ inbuffer_data[653];
assign xnor0[654] = 1'b1 ^~ inbuffer_data[654];
assign xnor0[655] = 1'b1 ^~ inbuffer_data[655];
assign xnor0[656] = 1'b1 ^~ inbuffer_data[656];
assign xnor0[657] = 1'b1 ^~ inbuffer_data[657];
assign xnor0[658] = 1'b1 ^~ inbuffer_data[658];
assign xnor0[659] = 1'b1 ^~ inbuffer_data[659];
assign xnor0[660] = 1'b0 ^~ inbuffer_data[660];
assign xnor0[661] = 1'b0 ^~ inbuffer_data[661];
assign xnor0[662] = 1'b0 ^~ inbuffer_data[662];
assign xnor0[663] = 1'b0 ^~ inbuffer_data[663];
assign xnor0[664] = 1'b0 ^~ inbuffer_data[664];
assign xnor0[665] = 1'b0 ^~ inbuffer_data[665];
assign xnor0[666] = 1'b0 ^~ inbuffer_data[666];
assign xnor0[667] = 1'b0 ^~ inbuffer_data[667];
assign xnor0[668] = 1'b1 ^~ inbuffer_data[668];
assign xnor0[669] = 1'b1 ^~ inbuffer_data[669];
assign xnor0[670] = 1'b0 ^~ inbuffer_data[670];
assign xnor0[671] = 1'b1 ^~ inbuffer_data[671];
assign xnor0[672] = 1'b1 ^~ inbuffer_data[672];
assign xnor0[673] = 1'b0 ^~ inbuffer_data[673];
assign xnor0[674] = 1'b1 ^~ inbuffer_data[674];
assign xnor0[675] = 1'b1 ^~ inbuffer_data[675];
assign xnor0[676] = 1'b1 ^~ inbuffer_data[676];
assign xnor0[677] = 1'b1 ^~ inbuffer_data[677];
assign xnor0[678] = 1'b0 ^~ inbuffer_data[678];
assign xnor0[679] = 1'b0 ^~ inbuffer_data[679];
assign xnor0[680] = 1'b0 ^~ inbuffer_data[680];
assign xnor0[681] = 1'b0 ^~ inbuffer_data[681];
assign xnor0[682] = 1'b1 ^~ inbuffer_data[682];
assign xnor0[683] = 1'b0 ^~ inbuffer_data[683];
assign xnor0[684] = 1'b1 ^~ inbuffer_data[684];
assign xnor0[685] = 1'b1 ^~ inbuffer_data[685];
assign xnor0[686] = 1'b1 ^~ inbuffer_data[686];
assign xnor0[687] = 1'b1 ^~ inbuffer_data[687];
assign xnor0[688] = 1'b1 ^~ inbuffer_data[688];
assign xnor0[689] = 1'b0 ^~ inbuffer_data[689];
assign xnor0[690] = 1'b0 ^~ inbuffer_data[690];
assign xnor0[691] = 1'b0 ^~ inbuffer_data[691];
assign xnor0[692] = 1'b0 ^~ inbuffer_data[692];
assign xnor0[693] = 1'b0 ^~ inbuffer_data[693];
assign xnor0[694] = 1'b1 ^~ inbuffer_data[694];
assign xnor0[695] = 1'b0 ^~ inbuffer_data[695];
assign xnor0[696] = 1'b0 ^~ inbuffer_data[696];
assign xnor0[697] = 1'b1 ^~ inbuffer_data[697];
assign xnor0[698] = 1'b0 ^~ inbuffer_data[698];
assign xnor0[699] = 1'b1 ^~ inbuffer_data[699];
assign xnor0[700] = 1'b1 ^~ inbuffer_data[700];
assign xnor0[701] = 1'b0 ^~ inbuffer_data[701];
assign xnor0[702] = 1'b0 ^~ inbuffer_data[702];
assign xnor0[703] = 1'b1 ^~ inbuffer_data[703];
assign xnor0[704] = 1'b1 ^~ inbuffer_data[704];
assign xnor0[705] = 1'b1 ^~ inbuffer_data[705];
assign xnor0[706] = 1'b0 ^~ inbuffer_data[706];
assign xnor0[707] = 1'b0 ^~ inbuffer_data[707];
assign xnor0[708] = 1'b0 ^~ inbuffer_data[708];
assign xnor0[709] = 1'b0 ^~ inbuffer_data[709];
assign xnor0[710] = 1'b0 ^~ inbuffer_data[710];
assign xnor0[711] = 1'b0 ^~ inbuffer_data[711];
assign xnor0[712] = 1'b0 ^~ inbuffer_data[712];
assign xnor0[713] = 1'b0 ^~ inbuffer_data[713];
assign xnor0[714] = 1'b0 ^~ inbuffer_data[714];
assign xnor0[715] = 1'b0 ^~ inbuffer_data[715];
assign xnor0[716] = 1'b0 ^~ inbuffer_data[716];
assign xnor0[717] = 1'b0 ^~ inbuffer_data[717];
assign xnor0[718] = 1'b0 ^~ inbuffer_data[718];
assign xnor0[719] = 1'b0 ^~ inbuffer_data[719];
assign xnor0[720] = 1'b0 ^~ inbuffer_data[720];
assign xnor0[721] = 1'b0 ^~ inbuffer_data[721];
assign xnor0[722] = 1'b0 ^~ inbuffer_data[722];
assign xnor0[723] = 1'b1 ^~ inbuffer_data[723];
assign xnor0[724] = 1'b1 ^~ inbuffer_data[724];
assign xnor0[725] = 1'b1 ^~ inbuffer_data[725];
assign xnor0[726] = 1'b1 ^~ inbuffer_data[726];
assign xnor0[727] = 1'b1 ^~ inbuffer_data[727];
assign xnor0[728] = 1'b0 ^~ inbuffer_data[728];
assign xnor0[729] = 1'b0 ^~ inbuffer_data[729];
assign xnor0[730] = 1'b1 ^~ inbuffer_data[730];
assign xnor0[731] = 1'b0 ^~ inbuffer_data[731];
assign xnor0[732] = 1'b1 ^~ inbuffer_data[732];
assign xnor0[733] = 1'b0 ^~ inbuffer_data[733];
assign xnor0[734] = 1'b0 ^~ inbuffer_data[734];
assign xnor0[735] = 1'b0 ^~ inbuffer_data[735];
assign xnor0[736] = 1'b0 ^~ inbuffer_data[736];
assign xnor0[737] = 1'b0 ^~ inbuffer_data[737];
assign xnor0[738] = 1'b0 ^~ inbuffer_data[738];
assign xnor0[739] = 1'b0 ^~ inbuffer_data[739];
assign xnor0[740] = 1'b0 ^~ inbuffer_data[740];
assign xnor0[741] = 1'b0 ^~ inbuffer_data[741];
assign xnor0[742] = 1'b0 ^~ inbuffer_data[742];
assign xnor0[743] = 1'b1 ^~ inbuffer_data[743];
assign xnor0[744] = 1'b1 ^~ inbuffer_data[744];
assign xnor0[745] = 1'b1 ^~ inbuffer_data[745];
assign xnor0[746] = 1'b1 ^~ inbuffer_data[746];
assign xnor0[747] = 1'b0 ^~ inbuffer_data[747];
assign xnor0[748] = 1'b0 ^~ inbuffer_data[748];
assign xnor0[749] = 1'b0 ^~ inbuffer_data[749];
assign xnor0[750] = 1'b1 ^~ inbuffer_data[750];
assign xnor0[751] = 1'b0 ^~ inbuffer_data[751];
assign xnor0[752] = 1'b1 ^~ inbuffer_data[752];
assign xnor0[753] = 1'b0 ^~ inbuffer_data[753];
assign xnor0[754] = 1'b0 ^~ inbuffer_data[754];
assign xnor0[755] = 1'b1 ^~ inbuffer_data[755];
assign xnor0[756] = 1'b0 ^~ inbuffer_data[756];
assign xnor0[757] = 1'b0 ^~ inbuffer_data[757];
assign xnor0[758] = 1'b0 ^~ inbuffer_data[758];
assign xnor0[759] = 1'b1 ^~ inbuffer_data[759];
assign xnor0[760] = 1'b0 ^~ inbuffer_data[760];
assign xnor0[761] = 1'b0 ^~ inbuffer_data[761];
assign xnor0[762] = 1'b0 ^~ inbuffer_data[762];
assign xnor0[763] = 1'b0 ^~ inbuffer_data[763];
assign xnor0[764] = 1'b1 ^~ inbuffer_data[764];
assign xnor0[765] = 1'b1 ^~ inbuffer_data[765];
assign xnor0[766] = 1'b0 ^~ inbuffer_data[766];
assign xnor0[767] = 1'b1 ^~ inbuffer_data[767];
assign xnor0[768] = 1'b0 ^~ inbuffer_data[768];
assign xnor0[769] = 1'b1 ^~ inbuffer_data[769];
assign xnor0[770] = 1'b1 ^~ inbuffer_data[770];
assign xnor0[771] = 1'b0 ^~ inbuffer_data[771];
assign xnor0[772] = 1'b1 ^~ inbuffer_data[772];
assign xnor0[773] = 1'b0 ^~ inbuffer_data[773];
assign xnor0[774] = 1'b1 ^~ inbuffer_data[774];
assign xnor0[775] = 1'b0 ^~ inbuffer_data[775];
assign xnor0[776] = 1'b1 ^~ inbuffer_data[776];
assign xnor0[777] = 1'b1 ^~ inbuffer_data[777];
assign xnor0[778] = 1'b0 ^~ inbuffer_data[778];
assign xnor0[779] = 1'b1 ^~ inbuffer_data[779];
assign xnor0[780] = 1'b0 ^~ inbuffer_data[780];
assign xnor0[781] = 1'b1 ^~ inbuffer_data[781];
assign xnor0[782] = 1'b1 ^~ inbuffer_data[782];
assign xnor0[783] = 1'b0 ^~ inbuffer_data[783];
assign xnor1[0] = 1'b0 ^~ inbuffer_data[0];
assign xnor1[1] = 1'b1 ^~ inbuffer_data[1];
assign xnor1[2] = 1'b1 ^~ inbuffer_data[2];
assign xnor1[3] = 1'b0 ^~ inbuffer_data[3];
assign xnor1[4] = 1'b0 ^~ inbuffer_data[4];
assign xnor1[5] = 1'b0 ^~ inbuffer_data[5];
assign xnor1[6] = 1'b1 ^~ inbuffer_data[6];
assign xnor1[7] = 1'b1 ^~ inbuffer_data[7];
assign xnor1[8] = 1'b1 ^~ inbuffer_data[8];
assign xnor1[9] = 1'b1 ^~ inbuffer_data[9];
assign xnor1[10] = 1'b1 ^~ inbuffer_data[10];
assign xnor1[11] = 1'b1 ^~ inbuffer_data[11];
assign xnor1[12] = 1'b0 ^~ inbuffer_data[12];
assign xnor1[13] = 1'b1 ^~ inbuffer_data[13];
assign xnor1[14] = 1'b0 ^~ inbuffer_data[14];
assign xnor1[15] = 1'b1 ^~ inbuffer_data[15];
assign xnor1[16] = 1'b1 ^~ inbuffer_data[16];
assign xnor1[17] = 1'b1 ^~ inbuffer_data[17];
assign xnor1[18] = 1'b1 ^~ inbuffer_data[18];
assign xnor1[19] = 1'b1 ^~ inbuffer_data[19];
assign xnor1[20] = 1'b0 ^~ inbuffer_data[20];
assign xnor1[21] = 1'b1 ^~ inbuffer_data[21];
assign xnor1[22] = 1'b1 ^~ inbuffer_data[22];
assign xnor1[23] = 1'b1 ^~ inbuffer_data[23];
assign xnor1[24] = 1'b0 ^~ inbuffer_data[24];
assign xnor1[25] = 1'b0 ^~ inbuffer_data[25];
assign xnor1[26] = 1'b1 ^~ inbuffer_data[26];
assign xnor1[27] = 1'b1 ^~ inbuffer_data[27];
assign xnor1[28] = 1'b1 ^~ inbuffer_data[28];
assign xnor1[29] = 1'b0 ^~ inbuffer_data[29];
assign xnor1[30] = 1'b1 ^~ inbuffer_data[30];
assign xnor1[31] = 1'b0 ^~ inbuffer_data[31];
assign xnor1[32] = 1'b0 ^~ inbuffer_data[32];
assign xnor1[33] = 1'b1 ^~ inbuffer_data[33];
assign xnor1[34] = 1'b0 ^~ inbuffer_data[34];
assign xnor1[35] = 1'b1 ^~ inbuffer_data[35];
assign xnor1[36] = 1'b1 ^~ inbuffer_data[36];
assign xnor1[37] = 1'b1 ^~ inbuffer_data[37];
assign xnor1[38] = 1'b1 ^~ inbuffer_data[38];
assign xnor1[39] = 1'b1 ^~ inbuffer_data[39];
assign xnor1[40] = 1'b0 ^~ inbuffer_data[40];
assign xnor1[41] = 1'b1 ^~ inbuffer_data[41];
assign xnor1[42] = 1'b1 ^~ inbuffer_data[42];
assign xnor1[43] = 1'b1 ^~ inbuffer_data[43];
assign xnor1[44] = 1'b1 ^~ inbuffer_data[44];
assign xnor1[45] = 1'b0 ^~ inbuffer_data[45];
assign xnor1[46] = 1'b1 ^~ inbuffer_data[46];
assign xnor1[47] = 1'b1 ^~ inbuffer_data[47];
assign xnor1[48] = 1'b1 ^~ inbuffer_data[48];
assign xnor1[49] = 1'b1 ^~ inbuffer_data[49];
assign xnor1[50] = 1'b0 ^~ inbuffer_data[50];
assign xnor1[51] = 1'b1 ^~ inbuffer_data[51];
assign xnor1[52] = 1'b0 ^~ inbuffer_data[52];
assign xnor1[53] = 1'b0 ^~ inbuffer_data[53];
assign xnor1[54] = 1'b1 ^~ inbuffer_data[54];
assign xnor1[55] = 1'b1 ^~ inbuffer_data[55];
assign xnor1[56] = 1'b0 ^~ inbuffer_data[56];
assign xnor1[57] = 1'b1 ^~ inbuffer_data[57];
assign xnor1[58] = 1'b0 ^~ inbuffer_data[58];
assign xnor1[59] = 1'b1 ^~ inbuffer_data[59];
assign xnor1[60] = 1'b1 ^~ inbuffer_data[60];
assign xnor1[61] = 1'b0 ^~ inbuffer_data[61];
assign xnor1[62] = 1'b0 ^~ inbuffer_data[62];
assign xnor1[63] = 1'b0 ^~ inbuffer_data[63];
assign xnor1[64] = 1'b0 ^~ inbuffer_data[64];
assign xnor1[65] = 1'b0 ^~ inbuffer_data[65];
assign xnor1[66] = 1'b0 ^~ inbuffer_data[66];
assign xnor1[67] = 1'b1 ^~ inbuffer_data[67];
assign xnor1[68] = 1'b1 ^~ inbuffer_data[68];
assign xnor1[69] = 1'b1 ^~ inbuffer_data[69];
assign xnor1[70] = 1'b0 ^~ inbuffer_data[70];
assign xnor1[71] = 1'b1 ^~ inbuffer_data[71];
assign xnor1[72] = 1'b1 ^~ inbuffer_data[72];
assign xnor1[73] = 1'b1 ^~ inbuffer_data[73];
assign xnor1[74] = 1'b0 ^~ inbuffer_data[74];
assign xnor1[75] = 1'b1 ^~ inbuffer_data[75];
assign xnor1[76] = 1'b1 ^~ inbuffer_data[76];
assign xnor1[77] = 1'b1 ^~ inbuffer_data[77];
assign xnor1[78] = 1'b1 ^~ inbuffer_data[78];
assign xnor1[79] = 1'b0 ^~ inbuffer_data[79];
assign xnor1[80] = 1'b0 ^~ inbuffer_data[80];
assign xnor1[81] = 1'b1 ^~ inbuffer_data[81];
assign xnor1[82] = 1'b0 ^~ inbuffer_data[82];
assign xnor1[83] = 1'b1 ^~ inbuffer_data[83];
assign xnor1[84] = 1'b0 ^~ inbuffer_data[84];
assign xnor1[85] = 1'b1 ^~ inbuffer_data[85];
assign xnor1[86] = 1'b1 ^~ inbuffer_data[86];
assign xnor1[87] = 1'b1 ^~ inbuffer_data[87];
assign xnor1[88] = 1'b0 ^~ inbuffer_data[88];
assign xnor1[89] = 1'b1 ^~ inbuffer_data[89];
assign xnor1[90] = 1'b0 ^~ inbuffer_data[90];
assign xnor1[91] = 1'b1 ^~ inbuffer_data[91];
assign xnor1[92] = 1'b1 ^~ inbuffer_data[92];
assign xnor1[93] = 1'b0 ^~ inbuffer_data[93];
assign xnor1[94] = 1'b1 ^~ inbuffer_data[94];
assign xnor1[95] = 1'b0 ^~ inbuffer_data[95];
assign xnor1[96] = 1'b1 ^~ inbuffer_data[96];
assign xnor1[97] = 1'b0 ^~ inbuffer_data[97];
assign xnor1[98] = 1'b1 ^~ inbuffer_data[98];
assign xnor1[99] = 1'b0 ^~ inbuffer_data[99];
assign xnor1[100] = 1'b0 ^~ inbuffer_data[100];
assign xnor1[101] = 1'b0 ^~ inbuffer_data[101];
assign xnor1[102] = 1'b0 ^~ inbuffer_data[102];
assign xnor1[103] = 1'b0 ^~ inbuffer_data[103];
assign xnor1[104] = 1'b0 ^~ inbuffer_data[104];
assign xnor1[105] = 1'b0 ^~ inbuffer_data[105];
assign xnor1[106] = 1'b1 ^~ inbuffer_data[106];
assign xnor1[107] = 1'b1 ^~ inbuffer_data[107];
assign xnor1[108] = 1'b0 ^~ inbuffer_data[108];
assign xnor1[109] = 1'b1 ^~ inbuffer_data[109];
assign xnor1[110] = 1'b0 ^~ inbuffer_data[110];
assign xnor1[111] = 1'b1 ^~ inbuffer_data[111];
assign xnor1[112] = 1'b0 ^~ inbuffer_data[112];
assign xnor1[113] = 1'b1 ^~ inbuffer_data[113];
assign xnor1[114] = 1'b0 ^~ inbuffer_data[114];
assign xnor1[115] = 1'b1 ^~ inbuffer_data[115];
assign xnor1[116] = 1'b0 ^~ inbuffer_data[116];
assign xnor1[117] = 1'b1 ^~ inbuffer_data[117];
assign xnor1[118] = 1'b1 ^~ inbuffer_data[118];
assign xnor1[119] = 1'b1 ^~ inbuffer_data[119];
assign xnor1[120] = 1'b0 ^~ inbuffer_data[120];
assign xnor1[121] = 1'b1 ^~ inbuffer_data[121];
assign xnor1[122] = 1'b0 ^~ inbuffer_data[122];
assign xnor1[123] = 1'b0 ^~ inbuffer_data[123];
assign xnor1[124] = 1'b0 ^~ inbuffer_data[124];
assign xnor1[125] = 1'b1 ^~ inbuffer_data[125];
assign xnor1[126] = 1'b0 ^~ inbuffer_data[126];
assign xnor1[127] = 1'b0 ^~ inbuffer_data[127];
assign xnor1[128] = 1'b1 ^~ inbuffer_data[128];
assign xnor1[129] = 1'b1 ^~ inbuffer_data[129];
assign xnor1[130] = 1'b1 ^~ inbuffer_data[130];
assign xnor1[131] = 1'b0 ^~ inbuffer_data[131];
assign xnor1[132] = 1'b1 ^~ inbuffer_data[132];
assign xnor1[133] = 1'b0 ^~ inbuffer_data[133];
assign xnor1[134] = 1'b0 ^~ inbuffer_data[134];
assign xnor1[135] = 1'b1 ^~ inbuffer_data[135];
assign xnor1[136] = 1'b0 ^~ inbuffer_data[136];
assign xnor1[137] = 1'b1 ^~ inbuffer_data[137];
assign xnor1[138] = 1'b1 ^~ inbuffer_data[138];
assign xnor1[139] = 1'b1 ^~ inbuffer_data[139];
assign xnor1[140] = 1'b0 ^~ inbuffer_data[140];
assign xnor1[141] = 1'b1 ^~ inbuffer_data[141];
assign xnor1[142] = 1'b0 ^~ inbuffer_data[142];
assign xnor1[143] = 1'b1 ^~ inbuffer_data[143];
assign xnor1[144] = 1'b1 ^~ inbuffer_data[144];
assign xnor1[145] = 1'b1 ^~ inbuffer_data[145];
assign xnor1[146] = 1'b1 ^~ inbuffer_data[146];
assign xnor1[147] = 1'b1 ^~ inbuffer_data[147];
assign xnor1[148] = 1'b0 ^~ inbuffer_data[148];
assign xnor1[149] = 1'b0 ^~ inbuffer_data[149];
assign xnor1[150] = 1'b0 ^~ inbuffer_data[150];
assign xnor1[151] = 1'b0 ^~ inbuffer_data[151];
assign xnor1[152] = 1'b1 ^~ inbuffer_data[152];
assign xnor1[153] = 1'b1 ^~ inbuffer_data[153];
assign xnor1[154] = 1'b0 ^~ inbuffer_data[154];
assign xnor1[155] = 1'b0 ^~ inbuffer_data[155];
assign xnor1[156] = 1'b1 ^~ inbuffer_data[156];
assign xnor1[157] = 1'b0 ^~ inbuffer_data[157];
assign xnor1[158] = 1'b0 ^~ inbuffer_data[158];
assign xnor1[159] = 1'b1 ^~ inbuffer_data[159];
assign xnor1[160] = 1'b0 ^~ inbuffer_data[160];
assign xnor1[161] = 1'b1 ^~ inbuffer_data[161];
assign xnor1[162] = 1'b1 ^~ inbuffer_data[162];
assign xnor1[163] = 1'b0 ^~ inbuffer_data[163];
assign xnor1[164] = 1'b1 ^~ inbuffer_data[164];
assign xnor1[165] = 1'b0 ^~ inbuffer_data[165];
assign xnor1[166] = 1'b1 ^~ inbuffer_data[166];
assign xnor1[167] = 1'b1 ^~ inbuffer_data[167];
assign xnor1[168] = 1'b0 ^~ inbuffer_data[168];
assign xnor1[169] = 1'b1 ^~ inbuffer_data[169];
assign xnor1[170] = 1'b1 ^~ inbuffer_data[170];
assign xnor1[171] = 1'b1 ^~ inbuffer_data[171];
assign xnor1[172] = 1'b1 ^~ inbuffer_data[172];
assign xnor1[173] = 1'b0 ^~ inbuffer_data[173];
assign xnor1[174] = 1'b1 ^~ inbuffer_data[174];
assign xnor1[175] = 1'b0 ^~ inbuffer_data[175];
assign xnor1[176] = 1'b0 ^~ inbuffer_data[176];
assign xnor1[177] = 1'b0 ^~ inbuffer_data[177];
assign xnor1[178] = 1'b0 ^~ inbuffer_data[178];
assign xnor1[179] = 1'b0 ^~ inbuffer_data[179];
assign xnor1[180] = 1'b0 ^~ inbuffer_data[180];
assign xnor1[181] = 1'b1 ^~ inbuffer_data[181];
assign xnor1[182] = 1'b0 ^~ inbuffer_data[182];
assign xnor1[183] = 1'b0 ^~ inbuffer_data[183];
assign xnor1[184] = 1'b0 ^~ inbuffer_data[184];
assign xnor1[185] = 1'b0 ^~ inbuffer_data[185];
assign xnor1[186] = 1'b0 ^~ inbuffer_data[186];
assign xnor1[187] = 1'b0 ^~ inbuffer_data[187];
assign xnor1[188] = 1'b1 ^~ inbuffer_data[188];
assign xnor1[189] = 1'b1 ^~ inbuffer_data[189];
assign xnor1[190] = 1'b0 ^~ inbuffer_data[190];
assign xnor1[191] = 1'b1 ^~ inbuffer_data[191];
assign xnor1[192] = 1'b0 ^~ inbuffer_data[192];
assign xnor1[193] = 1'b0 ^~ inbuffer_data[193];
assign xnor1[194] = 1'b0 ^~ inbuffer_data[194];
assign xnor1[195] = 1'b0 ^~ inbuffer_data[195];
assign xnor1[196] = 1'b1 ^~ inbuffer_data[196];
assign xnor1[197] = 1'b1 ^~ inbuffer_data[197];
assign xnor1[198] = 1'b1 ^~ inbuffer_data[198];
assign xnor1[199] = 1'b1 ^~ inbuffer_data[199];
assign xnor1[200] = 1'b1 ^~ inbuffer_data[200];
assign xnor1[201] = 1'b0 ^~ inbuffer_data[201];
assign xnor1[202] = 1'b0 ^~ inbuffer_data[202];
assign xnor1[203] = 1'b0 ^~ inbuffer_data[203];
assign xnor1[204] = 1'b0 ^~ inbuffer_data[204];
assign xnor1[205] = 1'b0 ^~ inbuffer_data[205];
assign xnor1[206] = 1'b0 ^~ inbuffer_data[206];
assign xnor1[207] = 1'b0 ^~ inbuffer_data[207];
assign xnor1[208] = 1'b0 ^~ inbuffer_data[208];
assign xnor1[209] = 1'b0 ^~ inbuffer_data[209];
assign xnor1[210] = 1'b0 ^~ inbuffer_data[210];
assign xnor1[211] = 1'b0 ^~ inbuffer_data[211];
assign xnor1[212] = 1'b0 ^~ inbuffer_data[212];
assign xnor1[213] = 1'b0 ^~ inbuffer_data[213];
assign xnor1[214] = 1'b0 ^~ inbuffer_data[214];
assign xnor1[215] = 1'b1 ^~ inbuffer_data[215];
assign xnor1[216] = 1'b1 ^~ inbuffer_data[216];
assign xnor1[217] = 1'b1 ^~ inbuffer_data[217];
assign xnor1[218] = 1'b0 ^~ inbuffer_data[218];
assign xnor1[219] = 1'b0 ^~ inbuffer_data[219];
assign xnor1[220] = 1'b0 ^~ inbuffer_data[220];
assign xnor1[221] = 1'b1 ^~ inbuffer_data[221];
assign xnor1[222] = 1'b1 ^~ inbuffer_data[222];
assign xnor1[223] = 1'b0 ^~ inbuffer_data[223];
assign xnor1[224] = 1'b1 ^~ inbuffer_data[224];
assign xnor1[225] = 1'b1 ^~ inbuffer_data[225];
assign xnor1[226] = 1'b1 ^~ inbuffer_data[226];
assign xnor1[227] = 1'b0 ^~ inbuffer_data[227];
assign xnor1[228] = 1'b1 ^~ inbuffer_data[228];
assign xnor1[229] = 1'b0 ^~ inbuffer_data[229];
assign xnor1[230] = 1'b0 ^~ inbuffer_data[230];
assign xnor1[231] = 1'b0 ^~ inbuffer_data[231];
assign xnor1[232] = 1'b0 ^~ inbuffer_data[232];
assign xnor1[233] = 1'b0 ^~ inbuffer_data[233];
assign xnor1[234] = 1'b0 ^~ inbuffer_data[234];
assign xnor1[235] = 1'b0 ^~ inbuffer_data[235];
assign xnor1[236] = 1'b1 ^~ inbuffer_data[236];
assign xnor1[237] = 1'b0 ^~ inbuffer_data[237];
assign xnor1[238] = 1'b1 ^~ inbuffer_data[238];
assign xnor1[239] = 1'b1 ^~ inbuffer_data[239];
assign xnor1[240] = 1'b0 ^~ inbuffer_data[240];
assign xnor1[241] = 1'b1 ^~ inbuffer_data[241];
assign xnor1[242] = 1'b1 ^~ inbuffer_data[242];
assign xnor1[243] = 1'b1 ^~ inbuffer_data[243];
assign xnor1[244] = 1'b0 ^~ inbuffer_data[244];
assign xnor1[245] = 1'b0 ^~ inbuffer_data[245];
assign xnor1[246] = 1'b0 ^~ inbuffer_data[246];
assign xnor1[247] = 1'b0 ^~ inbuffer_data[247];
assign xnor1[248] = 1'b0 ^~ inbuffer_data[248];
assign xnor1[249] = 1'b0 ^~ inbuffer_data[249];
assign xnor1[250] = 1'b0 ^~ inbuffer_data[250];
assign xnor1[251] = 1'b1 ^~ inbuffer_data[251];
assign xnor1[252] = 1'b1 ^~ inbuffer_data[252];
assign xnor1[253] = 1'b1 ^~ inbuffer_data[253];
assign xnor1[254] = 1'b1 ^~ inbuffer_data[254];
assign xnor1[255] = 1'b0 ^~ inbuffer_data[255];
assign xnor1[256] = 1'b0 ^~ inbuffer_data[256];
assign xnor1[257] = 1'b0 ^~ inbuffer_data[257];
assign xnor1[258] = 1'b0 ^~ inbuffer_data[258];
assign xnor1[259] = 1'b0 ^~ inbuffer_data[259];
assign xnor1[260] = 1'b0 ^~ inbuffer_data[260];
assign xnor1[261] = 1'b0 ^~ inbuffer_data[261];
assign xnor1[262] = 1'b0 ^~ inbuffer_data[262];
assign xnor1[263] = 1'b1 ^~ inbuffer_data[263];
assign xnor1[264] = 1'b1 ^~ inbuffer_data[264];
assign xnor1[265] = 1'b1 ^~ inbuffer_data[265];
assign xnor1[266] = 1'b1 ^~ inbuffer_data[266];
assign xnor1[267] = 1'b1 ^~ inbuffer_data[267];
assign xnor1[268] = 1'b1 ^~ inbuffer_data[268];
assign xnor1[269] = 1'b0 ^~ inbuffer_data[269];
assign xnor1[270] = 1'b1 ^~ inbuffer_data[270];
assign xnor1[271] = 1'b0 ^~ inbuffer_data[271];
assign xnor1[272] = 1'b0 ^~ inbuffer_data[272];
assign xnor1[273] = 1'b0 ^~ inbuffer_data[273];
assign xnor1[274] = 1'b0 ^~ inbuffer_data[274];
assign xnor1[275] = 1'b0 ^~ inbuffer_data[275];
assign xnor1[276] = 1'b0 ^~ inbuffer_data[276];
assign xnor1[277] = 1'b0 ^~ inbuffer_data[277];
assign xnor1[278] = 1'b0 ^~ inbuffer_data[278];
assign xnor1[279] = 1'b0 ^~ inbuffer_data[279];
assign xnor1[280] = 1'b1 ^~ inbuffer_data[280];
assign xnor1[281] = 1'b0 ^~ inbuffer_data[281];
assign xnor1[282] = 1'b0 ^~ inbuffer_data[282];
assign xnor1[283] = 1'b1 ^~ inbuffer_data[283];
assign xnor1[284] = 1'b1 ^~ inbuffer_data[284];
assign xnor1[285] = 1'b0 ^~ inbuffer_data[285];
assign xnor1[286] = 1'b0 ^~ inbuffer_data[286];
assign xnor1[287] = 1'b0 ^~ inbuffer_data[287];
assign xnor1[288] = 1'b0 ^~ inbuffer_data[288];
assign xnor1[289] = 1'b0 ^~ inbuffer_data[289];
assign xnor1[290] = 1'b1 ^~ inbuffer_data[290];
assign xnor1[291] = 1'b0 ^~ inbuffer_data[291];
assign xnor1[292] = 1'b0 ^~ inbuffer_data[292];
assign xnor1[293] = 1'b1 ^~ inbuffer_data[293];
assign xnor1[294] = 1'b1 ^~ inbuffer_data[294];
assign xnor1[295] = 1'b1 ^~ inbuffer_data[295];
assign xnor1[296] = 1'b1 ^~ inbuffer_data[296];
assign xnor1[297] = 1'b1 ^~ inbuffer_data[297];
assign xnor1[298] = 1'b0 ^~ inbuffer_data[298];
assign xnor1[299] = 1'b0 ^~ inbuffer_data[299];
assign xnor1[300] = 1'b0 ^~ inbuffer_data[300];
assign xnor1[301] = 1'b0 ^~ inbuffer_data[301];
assign xnor1[302] = 1'b0 ^~ inbuffer_data[302];
assign xnor1[303] = 1'b0 ^~ inbuffer_data[303];
assign xnor1[304] = 1'b0 ^~ inbuffer_data[304];
assign xnor1[305] = 1'b0 ^~ inbuffer_data[305];
assign xnor1[306] = 1'b0 ^~ inbuffer_data[306];
assign xnor1[307] = 1'b0 ^~ inbuffer_data[307];
assign xnor1[308] = 1'b1 ^~ inbuffer_data[308];
assign xnor1[309] = 1'b1 ^~ inbuffer_data[309];
assign xnor1[310] = 1'b1 ^~ inbuffer_data[310];
assign xnor1[311] = 1'b1 ^~ inbuffer_data[311];
assign xnor1[312] = 1'b1 ^~ inbuffer_data[312];
assign xnor1[313] = 1'b0 ^~ inbuffer_data[313];
assign xnor1[314] = 1'b1 ^~ inbuffer_data[314];
assign xnor1[315] = 1'b0 ^~ inbuffer_data[315];
assign xnor1[316] = 1'b1 ^~ inbuffer_data[316];
assign xnor1[317] = 1'b0 ^~ inbuffer_data[317];
assign xnor1[318] = 1'b1 ^~ inbuffer_data[318];
assign xnor1[319] = 1'b0 ^~ inbuffer_data[319];
assign xnor1[320] = 1'b0 ^~ inbuffer_data[320];
assign xnor1[321] = 1'b1 ^~ inbuffer_data[321];
assign xnor1[322] = 1'b1 ^~ inbuffer_data[322];
assign xnor1[323] = 1'b1 ^~ inbuffer_data[323];
assign xnor1[324] = 1'b1 ^~ inbuffer_data[324];
assign xnor1[325] = 1'b0 ^~ inbuffer_data[325];
assign xnor1[326] = 1'b1 ^~ inbuffer_data[326];
assign xnor1[327] = 1'b0 ^~ inbuffer_data[327];
assign xnor1[328] = 1'b0 ^~ inbuffer_data[328];
assign xnor1[329] = 1'b0 ^~ inbuffer_data[329];
assign xnor1[330] = 1'b0 ^~ inbuffer_data[330];
assign xnor1[331] = 1'b0 ^~ inbuffer_data[331];
assign xnor1[332] = 1'b0 ^~ inbuffer_data[332];
assign xnor1[333] = 1'b0 ^~ inbuffer_data[333];
assign xnor1[334] = 1'b0 ^~ inbuffer_data[334];
assign xnor1[335] = 1'b0 ^~ inbuffer_data[335];
assign xnor1[336] = 1'b0 ^~ inbuffer_data[336];
assign xnor1[337] = 1'b0 ^~ inbuffer_data[337];
assign xnor1[338] = 1'b1 ^~ inbuffer_data[338];
assign xnor1[339] = 1'b1 ^~ inbuffer_data[339];
assign xnor1[340] = 1'b1 ^~ inbuffer_data[340];
assign xnor1[341] = 1'b0 ^~ inbuffer_data[341];
assign xnor1[342] = 1'b0 ^~ inbuffer_data[342];
assign xnor1[343] = 1'b0 ^~ inbuffer_data[343];
assign xnor1[344] = 1'b0 ^~ inbuffer_data[344];
assign xnor1[345] = 1'b1 ^~ inbuffer_data[345];
assign xnor1[346] = 1'b0 ^~ inbuffer_data[346];
assign xnor1[347] = 1'b0 ^~ inbuffer_data[347];
assign xnor1[348] = 1'b0 ^~ inbuffer_data[348];
assign xnor1[349] = 1'b1 ^~ inbuffer_data[349];
assign xnor1[350] = 1'b1 ^~ inbuffer_data[350];
assign xnor1[351] = 1'b1 ^~ inbuffer_data[351];
assign xnor1[352] = 1'b1 ^~ inbuffer_data[352];
assign xnor1[353] = 1'b0 ^~ inbuffer_data[353];
assign xnor1[354] = 1'b0 ^~ inbuffer_data[354];
assign xnor1[355] = 1'b0 ^~ inbuffer_data[355];
assign xnor1[356] = 1'b0 ^~ inbuffer_data[356];
assign xnor1[357] = 1'b1 ^~ inbuffer_data[357];
assign xnor1[358] = 1'b0 ^~ inbuffer_data[358];
assign xnor1[359] = 1'b0 ^~ inbuffer_data[359];
assign xnor1[360] = 1'b0 ^~ inbuffer_data[360];
assign xnor1[361] = 1'b1 ^~ inbuffer_data[361];
assign xnor1[362] = 1'b1 ^~ inbuffer_data[362];
assign xnor1[363] = 1'b1 ^~ inbuffer_data[363];
assign xnor1[364] = 1'b1 ^~ inbuffer_data[364];
assign xnor1[365] = 1'b1 ^~ inbuffer_data[365];
assign xnor1[366] = 1'b1 ^~ inbuffer_data[366];
assign xnor1[367] = 1'b1 ^~ inbuffer_data[367];
assign xnor1[368] = 1'b0 ^~ inbuffer_data[368];
assign xnor1[369] = 1'b1 ^~ inbuffer_data[369];
assign xnor1[370] = 1'b1 ^~ inbuffer_data[370];
assign xnor1[371] = 1'b0 ^~ inbuffer_data[371];
assign xnor1[372] = 1'b1 ^~ inbuffer_data[372];
assign xnor1[373] = 1'b0 ^~ inbuffer_data[373];
assign xnor1[374] = 1'b0 ^~ inbuffer_data[374];
assign xnor1[375] = 1'b0 ^~ inbuffer_data[375];
assign xnor1[376] = 1'b0 ^~ inbuffer_data[376];
assign xnor1[377] = 1'b1 ^~ inbuffer_data[377];
assign xnor1[378] = 1'b1 ^~ inbuffer_data[378];
assign xnor1[379] = 1'b1 ^~ inbuffer_data[379];
assign xnor1[380] = 1'b0 ^~ inbuffer_data[380];
assign xnor1[381] = 1'b0 ^~ inbuffer_data[381];
assign xnor1[382] = 1'b0 ^~ inbuffer_data[382];
assign xnor1[383] = 1'b0 ^~ inbuffer_data[383];
assign xnor1[384] = 1'b0 ^~ inbuffer_data[384];
assign xnor1[385] = 1'b0 ^~ inbuffer_data[385];
assign xnor1[386] = 1'b0 ^~ inbuffer_data[386];
assign xnor1[387] = 1'b1 ^~ inbuffer_data[387];
assign xnor1[388] = 1'b1 ^~ inbuffer_data[388];
assign xnor1[389] = 1'b0 ^~ inbuffer_data[389];
assign xnor1[390] = 1'b1 ^~ inbuffer_data[390];
assign xnor1[391] = 1'b1 ^~ inbuffer_data[391];
assign xnor1[392] = 1'b1 ^~ inbuffer_data[392];
assign xnor1[393] = 1'b0 ^~ inbuffer_data[393];
assign xnor1[394] = 1'b0 ^~ inbuffer_data[394];
assign xnor1[395] = 1'b0 ^~ inbuffer_data[395];
assign xnor1[396] = 1'b1 ^~ inbuffer_data[396];
assign xnor1[397] = 1'b1 ^~ inbuffer_data[397];
assign xnor1[398] = 1'b0 ^~ inbuffer_data[398];
assign xnor1[399] = 1'b0 ^~ inbuffer_data[399];
assign xnor1[400] = 1'b0 ^~ inbuffer_data[400];
assign xnor1[401] = 1'b0 ^~ inbuffer_data[401];
assign xnor1[402] = 1'b0 ^~ inbuffer_data[402];
assign xnor1[403] = 1'b0 ^~ inbuffer_data[403];
assign xnor1[404] = 1'b1 ^~ inbuffer_data[404];
assign xnor1[405] = 1'b1 ^~ inbuffer_data[405];
assign xnor1[406] = 1'b1 ^~ inbuffer_data[406];
assign xnor1[407] = 1'b1 ^~ inbuffer_data[407];
assign xnor1[408] = 1'b1 ^~ inbuffer_data[408];
assign xnor1[409] = 1'b0 ^~ inbuffer_data[409];
assign xnor1[410] = 1'b0 ^~ inbuffer_data[410];
assign xnor1[411] = 1'b0 ^~ inbuffer_data[411];
assign xnor1[412] = 1'b0 ^~ inbuffer_data[412];
assign xnor1[413] = 1'b1 ^~ inbuffer_data[413];
assign xnor1[414] = 1'b1 ^~ inbuffer_data[414];
assign xnor1[415] = 1'b1 ^~ inbuffer_data[415];
assign xnor1[416] = 1'b0 ^~ inbuffer_data[416];
assign xnor1[417] = 1'b1 ^~ inbuffer_data[417];
assign xnor1[418] = 1'b1 ^~ inbuffer_data[418];
assign xnor1[419] = 1'b0 ^~ inbuffer_data[419];
assign xnor1[420] = 1'b1 ^~ inbuffer_data[420];
assign xnor1[421] = 1'b1 ^~ inbuffer_data[421];
assign xnor1[422] = 1'b1 ^~ inbuffer_data[422];
assign xnor1[423] = 1'b1 ^~ inbuffer_data[423];
assign xnor1[424] = 1'b0 ^~ inbuffer_data[424];
assign xnor1[425] = 1'b0 ^~ inbuffer_data[425];
assign xnor1[426] = 1'b0 ^~ inbuffer_data[426];
assign xnor1[427] = 1'b0 ^~ inbuffer_data[427];
assign xnor1[428] = 1'b1 ^~ inbuffer_data[428];
assign xnor1[429] = 1'b0 ^~ inbuffer_data[429];
assign xnor1[430] = 1'b0 ^~ inbuffer_data[430];
assign xnor1[431] = 1'b0 ^~ inbuffer_data[431];
assign xnor1[432] = 1'b0 ^~ inbuffer_data[432];
assign xnor1[433] = 1'b1 ^~ inbuffer_data[433];
assign xnor1[434] = 1'b1 ^~ inbuffer_data[434];
assign xnor1[435] = 1'b1 ^~ inbuffer_data[435];
assign xnor1[436] = 1'b0 ^~ inbuffer_data[436];
assign xnor1[437] = 1'b0 ^~ inbuffer_data[437];
assign xnor1[438] = 1'b0 ^~ inbuffer_data[438];
assign xnor1[439] = 1'b0 ^~ inbuffer_data[439];
assign xnor1[440] = 1'b0 ^~ inbuffer_data[440];
assign xnor1[441] = 1'b0 ^~ inbuffer_data[441];
assign xnor1[442] = 1'b0 ^~ inbuffer_data[442];
assign xnor1[443] = 1'b1 ^~ inbuffer_data[443];
assign xnor1[444] = 1'b0 ^~ inbuffer_data[444];
assign xnor1[445] = 1'b0 ^~ inbuffer_data[445];
assign xnor1[446] = 1'b0 ^~ inbuffer_data[446];
assign xnor1[447] = 1'b0 ^~ inbuffer_data[447];
assign xnor1[448] = 1'b1 ^~ inbuffer_data[448];
assign xnor1[449] = 1'b1 ^~ inbuffer_data[449];
assign xnor1[450] = 1'b1 ^~ inbuffer_data[450];
assign xnor1[451] = 1'b0 ^~ inbuffer_data[451];
assign xnor1[452] = 1'b1 ^~ inbuffer_data[452];
assign xnor1[453] = 1'b0 ^~ inbuffer_data[453];
assign xnor1[454] = 1'b0 ^~ inbuffer_data[454];
assign xnor1[455] = 1'b0 ^~ inbuffer_data[455];
assign xnor1[456] = 1'b0 ^~ inbuffer_data[456];
assign xnor1[457] = 1'b0 ^~ inbuffer_data[457];
assign xnor1[458] = 1'b0 ^~ inbuffer_data[458];
assign xnor1[459] = 1'b0 ^~ inbuffer_data[459];
assign xnor1[460] = 1'b0 ^~ inbuffer_data[460];
assign xnor1[461] = 1'b1 ^~ inbuffer_data[461];
assign xnor1[462] = 1'b1 ^~ inbuffer_data[462];
assign xnor1[463] = 1'b1 ^~ inbuffer_data[463];
assign xnor1[464] = 1'b0 ^~ inbuffer_data[464];
assign xnor1[465] = 1'b0 ^~ inbuffer_data[465];
assign xnor1[466] = 1'b0 ^~ inbuffer_data[466];
assign xnor1[467] = 1'b0 ^~ inbuffer_data[467];
assign xnor1[468] = 1'b0 ^~ inbuffer_data[468];
assign xnor1[469] = 1'b0 ^~ inbuffer_data[469];
assign xnor1[470] = 1'b0 ^~ inbuffer_data[470];
assign xnor1[471] = 1'b0 ^~ inbuffer_data[471];
assign xnor1[472] = 1'b1 ^~ inbuffer_data[472];
assign xnor1[473] = 1'b0 ^~ inbuffer_data[473];
assign xnor1[474] = 1'b1 ^~ inbuffer_data[474];
assign xnor1[475] = 1'b1 ^~ inbuffer_data[475];
assign xnor1[476] = 1'b0 ^~ inbuffer_data[476];
assign xnor1[477] = 1'b0 ^~ inbuffer_data[477];
assign xnor1[478] = 1'b1 ^~ inbuffer_data[478];
assign xnor1[479] = 1'b0 ^~ inbuffer_data[479];
assign xnor1[480] = 1'b1 ^~ inbuffer_data[480];
assign xnor1[481] = 1'b0 ^~ inbuffer_data[481];
assign xnor1[482] = 1'b0 ^~ inbuffer_data[482];
assign xnor1[483] = 1'b0 ^~ inbuffer_data[483];
assign xnor1[484] = 1'b0 ^~ inbuffer_data[484];
assign xnor1[485] = 1'b1 ^~ inbuffer_data[485];
assign xnor1[486] = 1'b1 ^~ inbuffer_data[486];
assign xnor1[487] = 1'b0 ^~ inbuffer_data[487];
assign xnor1[488] = 1'b1 ^~ inbuffer_data[488];
assign xnor1[489] = 1'b1 ^~ inbuffer_data[489];
assign xnor1[490] = 1'b1 ^~ inbuffer_data[490];
assign xnor1[491] = 1'b1 ^~ inbuffer_data[491];
assign xnor1[492] = 1'b0 ^~ inbuffer_data[492];
assign xnor1[493] = 1'b0 ^~ inbuffer_data[493];
assign xnor1[494] = 1'b0 ^~ inbuffer_data[494];
assign xnor1[495] = 1'b0 ^~ inbuffer_data[495];
assign xnor1[496] = 1'b0 ^~ inbuffer_data[496];
assign xnor1[497] = 1'b0 ^~ inbuffer_data[497];
assign xnor1[498] = 1'b0 ^~ inbuffer_data[498];
assign xnor1[499] = 1'b1 ^~ inbuffer_data[499];
assign xnor1[500] = 1'b0 ^~ inbuffer_data[500];
assign xnor1[501] = 1'b0 ^~ inbuffer_data[501];
assign xnor1[502] = 1'b1 ^~ inbuffer_data[502];
assign xnor1[503] = 1'b1 ^~ inbuffer_data[503];
assign xnor1[504] = 1'b1 ^~ inbuffer_data[504];
assign xnor1[505] = 1'b0 ^~ inbuffer_data[505];
assign xnor1[506] = 1'b0 ^~ inbuffer_data[506];
assign xnor1[507] = 1'b1 ^~ inbuffer_data[507];
assign xnor1[508] = 1'b0 ^~ inbuffer_data[508];
assign xnor1[509] = 1'b0 ^~ inbuffer_data[509];
assign xnor1[510] = 1'b0 ^~ inbuffer_data[510];
assign xnor1[511] = 1'b0 ^~ inbuffer_data[511];
assign xnor1[512] = 1'b1 ^~ inbuffer_data[512];
assign xnor1[513] = 1'b0 ^~ inbuffer_data[513];
assign xnor1[514] = 1'b0 ^~ inbuffer_data[514];
assign xnor1[515] = 1'b1 ^~ inbuffer_data[515];
assign xnor1[516] = 1'b1 ^~ inbuffer_data[516];
assign xnor1[517] = 1'b1 ^~ inbuffer_data[517];
assign xnor1[518] = 1'b1 ^~ inbuffer_data[518];
assign xnor1[519] = 1'b0 ^~ inbuffer_data[519];
assign xnor1[520] = 1'b0 ^~ inbuffer_data[520];
assign xnor1[521] = 1'b0 ^~ inbuffer_data[521];
assign xnor1[522] = 1'b0 ^~ inbuffer_data[522];
assign xnor1[523] = 1'b1 ^~ inbuffer_data[523];
assign xnor1[524] = 1'b0 ^~ inbuffer_data[524];
assign xnor1[525] = 1'b1 ^~ inbuffer_data[525];
assign xnor1[526] = 1'b0 ^~ inbuffer_data[526];
assign xnor1[527] = 1'b0 ^~ inbuffer_data[527];
assign xnor1[528] = 1'b0 ^~ inbuffer_data[528];
assign xnor1[529] = 1'b1 ^~ inbuffer_data[529];
assign xnor1[530] = 1'b0 ^~ inbuffer_data[530];
assign xnor1[531] = 1'b1 ^~ inbuffer_data[531];
assign xnor1[532] = 1'b1 ^~ inbuffer_data[532];
assign xnor1[533] = 1'b1 ^~ inbuffer_data[533];
assign xnor1[534] = 1'b0 ^~ inbuffer_data[534];
assign xnor1[535] = 1'b0 ^~ inbuffer_data[535];
assign xnor1[536] = 1'b1 ^~ inbuffer_data[536];
assign xnor1[537] = 1'b0 ^~ inbuffer_data[537];
assign xnor1[538] = 1'b0 ^~ inbuffer_data[538];
assign xnor1[539] = 1'b0 ^~ inbuffer_data[539];
assign xnor1[540] = 1'b0 ^~ inbuffer_data[540];
assign xnor1[541] = 1'b1 ^~ inbuffer_data[541];
assign xnor1[542] = 1'b0 ^~ inbuffer_data[542];
assign xnor1[543] = 1'b1 ^~ inbuffer_data[543];
assign xnor1[544] = 1'b0 ^~ inbuffer_data[544];
assign xnor1[545] = 1'b1 ^~ inbuffer_data[545];
assign xnor1[546] = 1'b1 ^~ inbuffer_data[546];
assign xnor1[547] = 1'b1 ^~ inbuffer_data[547];
assign xnor1[548] = 1'b1 ^~ inbuffer_data[548];
assign xnor1[549] = 1'b0 ^~ inbuffer_data[549];
assign xnor1[550] = 1'b1 ^~ inbuffer_data[550];
assign xnor1[551] = 1'b0 ^~ inbuffer_data[551];
assign xnor1[552] = 1'b1 ^~ inbuffer_data[552];
assign xnor1[553] = 1'b0 ^~ inbuffer_data[553];
assign xnor1[554] = 1'b0 ^~ inbuffer_data[554];
assign xnor1[555] = 1'b0 ^~ inbuffer_data[555];
assign xnor1[556] = 1'b0 ^~ inbuffer_data[556];
assign xnor1[557] = 1'b1 ^~ inbuffer_data[557];
assign xnor1[558] = 1'b1 ^~ inbuffer_data[558];
assign xnor1[559] = 1'b1 ^~ inbuffer_data[559];
assign xnor1[560] = 1'b1 ^~ inbuffer_data[560];
assign xnor1[561] = 1'b1 ^~ inbuffer_data[561];
assign xnor1[562] = 1'b1 ^~ inbuffer_data[562];
assign xnor1[563] = 1'b0 ^~ inbuffer_data[563];
assign xnor1[564] = 1'b1 ^~ inbuffer_data[564];
assign xnor1[565] = 1'b0 ^~ inbuffer_data[565];
assign xnor1[566] = 1'b1 ^~ inbuffer_data[566];
assign xnor1[567] = 1'b0 ^~ inbuffer_data[567];
assign xnor1[568] = 1'b1 ^~ inbuffer_data[568];
assign xnor1[569] = 1'b1 ^~ inbuffer_data[569];
assign xnor1[570] = 1'b1 ^~ inbuffer_data[570];
assign xnor1[571] = 1'b1 ^~ inbuffer_data[571];
assign xnor1[572] = 1'b1 ^~ inbuffer_data[572];
assign xnor1[573] = 1'b1 ^~ inbuffer_data[573];
assign xnor1[574] = 1'b0 ^~ inbuffer_data[574];
assign xnor1[575] = 1'b0 ^~ inbuffer_data[575];
assign xnor1[576] = 1'b1 ^~ inbuffer_data[576];
assign xnor1[577] = 1'b1 ^~ inbuffer_data[577];
assign xnor1[578] = 1'b0 ^~ inbuffer_data[578];
assign xnor1[579] = 1'b1 ^~ inbuffer_data[579];
assign xnor1[580] = 1'b1 ^~ inbuffer_data[580];
assign xnor1[581] = 1'b1 ^~ inbuffer_data[581];
assign xnor1[582] = 1'b0 ^~ inbuffer_data[582];
assign xnor1[583] = 1'b0 ^~ inbuffer_data[583];
assign xnor1[584] = 1'b1 ^~ inbuffer_data[584];
assign xnor1[585] = 1'b1 ^~ inbuffer_data[585];
assign xnor1[586] = 1'b0 ^~ inbuffer_data[586];
assign xnor1[587] = 1'b0 ^~ inbuffer_data[587];
assign xnor1[588] = 1'b1 ^~ inbuffer_data[588];
assign xnor1[589] = 1'b1 ^~ inbuffer_data[589];
assign xnor1[590] = 1'b0 ^~ inbuffer_data[590];
assign xnor1[591] = 1'b1 ^~ inbuffer_data[591];
assign xnor1[592] = 1'b1 ^~ inbuffer_data[592];
assign xnor1[593] = 1'b1 ^~ inbuffer_data[593];
assign xnor1[594] = 1'b1 ^~ inbuffer_data[594];
assign xnor1[595] = 1'b1 ^~ inbuffer_data[595];
assign xnor1[596] = 1'b1 ^~ inbuffer_data[596];
assign xnor1[597] = 1'b1 ^~ inbuffer_data[597];
assign xnor1[598] = 1'b1 ^~ inbuffer_data[598];
assign xnor1[599] = 1'b0 ^~ inbuffer_data[599];
assign xnor1[600] = 1'b0 ^~ inbuffer_data[600];
assign xnor1[601] = 1'b0 ^~ inbuffer_data[601];
assign xnor1[602] = 1'b0 ^~ inbuffer_data[602];
assign xnor1[603] = 1'b1 ^~ inbuffer_data[603];
assign xnor1[604] = 1'b1 ^~ inbuffer_data[604];
assign xnor1[605] = 1'b1 ^~ inbuffer_data[605];
assign xnor1[606] = 1'b1 ^~ inbuffer_data[606];
assign xnor1[607] = 1'b1 ^~ inbuffer_data[607];
assign xnor1[608] = 1'b1 ^~ inbuffer_data[608];
assign xnor1[609] = 1'b0 ^~ inbuffer_data[609];
assign xnor1[610] = 1'b0 ^~ inbuffer_data[610];
assign xnor1[611] = 1'b1 ^~ inbuffer_data[611];
assign xnor1[612] = 1'b1 ^~ inbuffer_data[612];
assign xnor1[613] = 1'b1 ^~ inbuffer_data[613];
assign xnor1[614] = 1'b0 ^~ inbuffer_data[614];
assign xnor1[615] = 1'b1 ^~ inbuffer_data[615];
assign xnor1[616] = 1'b1 ^~ inbuffer_data[616];
assign xnor1[617] = 1'b0 ^~ inbuffer_data[617];
assign xnor1[618] = 1'b0 ^~ inbuffer_data[618];
assign xnor1[619] = 1'b1 ^~ inbuffer_data[619];
assign xnor1[620] = 1'b0 ^~ inbuffer_data[620];
assign xnor1[621] = 1'b1 ^~ inbuffer_data[621];
assign xnor1[622] = 1'b1 ^~ inbuffer_data[622];
assign xnor1[623] = 1'b1 ^~ inbuffer_data[623];
assign xnor1[624] = 1'b0 ^~ inbuffer_data[624];
assign xnor1[625] = 1'b1 ^~ inbuffer_data[625];
assign xnor1[626] = 1'b1 ^~ inbuffer_data[626];
assign xnor1[627] = 1'b0 ^~ inbuffer_data[627];
assign xnor1[628] = 1'b0 ^~ inbuffer_data[628];
assign xnor1[629] = 1'b0 ^~ inbuffer_data[629];
assign xnor1[630] = 1'b0 ^~ inbuffer_data[630];
assign xnor1[631] = 1'b0 ^~ inbuffer_data[631];
assign xnor1[632] = 1'b1 ^~ inbuffer_data[632];
assign xnor1[633] = 1'b1 ^~ inbuffer_data[633];
assign xnor1[634] = 1'b1 ^~ inbuffer_data[634];
assign xnor1[635] = 1'b1 ^~ inbuffer_data[635];
assign xnor1[636] = 1'b1 ^~ inbuffer_data[636];
assign xnor1[637] = 1'b1 ^~ inbuffer_data[637];
assign xnor1[638] = 1'b0 ^~ inbuffer_data[638];
assign xnor1[639] = 1'b1 ^~ inbuffer_data[639];
assign xnor1[640] = 1'b0 ^~ inbuffer_data[640];
assign xnor1[641] = 1'b1 ^~ inbuffer_data[641];
assign xnor1[642] = 1'b1 ^~ inbuffer_data[642];
assign xnor1[643] = 1'b0 ^~ inbuffer_data[643];
assign xnor1[644] = 1'b0 ^~ inbuffer_data[644];
assign xnor1[645] = 1'b0 ^~ inbuffer_data[645];
assign xnor1[646] = 1'b0 ^~ inbuffer_data[646];
assign xnor1[647] = 1'b1 ^~ inbuffer_data[647];
assign xnor1[648] = 1'b1 ^~ inbuffer_data[648];
assign xnor1[649] = 1'b1 ^~ inbuffer_data[649];
assign xnor1[650] = 1'b1 ^~ inbuffer_data[650];
assign xnor1[651] = 1'b1 ^~ inbuffer_data[651];
assign xnor1[652] = 1'b1 ^~ inbuffer_data[652];
assign xnor1[653] = 1'b1 ^~ inbuffer_data[653];
assign xnor1[654] = 1'b0 ^~ inbuffer_data[654];
assign xnor1[655] = 1'b1 ^~ inbuffer_data[655];
assign xnor1[656] = 1'b0 ^~ inbuffer_data[656];
assign xnor1[657] = 1'b1 ^~ inbuffer_data[657];
assign xnor1[658] = 1'b0 ^~ inbuffer_data[658];
assign xnor1[659] = 1'b1 ^~ inbuffer_data[659];
assign xnor1[660] = 1'b1 ^~ inbuffer_data[660];
assign xnor1[661] = 1'b1 ^~ inbuffer_data[661];
assign xnor1[662] = 1'b1 ^~ inbuffer_data[662];
assign xnor1[663] = 1'b1 ^~ inbuffer_data[663];
assign xnor1[664] = 1'b0 ^~ inbuffer_data[664];
assign xnor1[665] = 1'b0 ^~ inbuffer_data[665];
assign xnor1[666] = 1'b0 ^~ inbuffer_data[666];
assign xnor1[667] = 1'b0 ^~ inbuffer_data[667];
assign xnor1[668] = 1'b0 ^~ inbuffer_data[668];
assign xnor1[669] = 1'b1 ^~ inbuffer_data[669];
assign xnor1[670] = 1'b0 ^~ inbuffer_data[670];
assign xnor1[671] = 1'b1 ^~ inbuffer_data[671];
assign xnor1[672] = 1'b0 ^~ inbuffer_data[672];
assign xnor1[673] = 1'b1 ^~ inbuffer_data[673];
assign xnor1[674] = 1'b1 ^~ inbuffer_data[674];
assign xnor1[675] = 1'b1 ^~ inbuffer_data[675];
assign xnor1[676] = 1'b1 ^~ inbuffer_data[676];
assign xnor1[677] = 1'b1 ^~ inbuffer_data[677];
assign xnor1[678] = 1'b0 ^~ inbuffer_data[678];
assign xnor1[679] = 1'b0 ^~ inbuffer_data[679];
assign xnor1[680] = 1'b0 ^~ inbuffer_data[680];
assign xnor1[681] = 1'b1 ^~ inbuffer_data[681];
assign xnor1[682] = 1'b0 ^~ inbuffer_data[682];
assign xnor1[683] = 1'b0 ^~ inbuffer_data[683];
assign xnor1[684] = 1'b0 ^~ inbuffer_data[684];
assign xnor1[685] = 1'b0 ^~ inbuffer_data[685];
assign xnor1[686] = 1'b0 ^~ inbuffer_data[686];
assign xnor1[687] = 1'b0 ^~ inbuffer_data[687];
assign xnor1[688] = 1'b0 ^~ inbuffer_data[688];
assign xnor1[689] = 1'b0 ^~ inbuffer_data[689];
assign xnor1[690] = 1'b1 ^~ inbuffer_data[690];
assign xnor1[691] = 1'b1 ^~ inbuffer_data[691];
assign xnor1[692] = 1'b0 ^~ inbuffer_data[692];
assign xnor1[693] = 1'b0 ^~ inbuffer_data[693];
assign xnor1[694] = 1'b1 ^~ inbuffer_data[694];
assign xnor1[695] = 1'b1 ^~ inbuffer_data[695];
assign xnor1[696] = 1'b1 ^~ inbuffer_data[696];
assign xnor1[697] = 1'b1 ^~ inbuffer_data[697];
assign xnor1[698] = 1'b1 ^~ inbuffer_data[698];
assign xnor1[699] = 1'b0 ^~ inbuffer_data[699];
assign xnor1[700] = 1'b1 ^~ inbuffer_data[700];
assign xnor1[701] = 1'b1 ^~ inbuffer_data[701];
assign xnor1[702] = 1'b1 ^~ inbuffer_data[702];
assign xnor1[703] = 1'b1 ^~ inbuffer_data[703];
assign xnor1[704] = 1'b1 ^~ inbuffer_data[704];
assign xnor1[705] = 1'b0 ^~ inbuffer_data[705];
assign xnor1[706] = 1'b0 ^~ inbuffer_data[706];
assign xnor1[707] = 1'b0 ^~ inbuffer_data[707];
assign xnor1[708] = 1'b0 ^~ inbuffer_data[708];
assign xnor1[709] = 1'b0 ^~ inbuffer_data[709];
assign xnor1[710] = 1'b0 ^~ inbuffer_data[710];
assign xnor1[711] = 1'b0 ^~ inbuffer_data[711];
assign xnor1[712] = 1'b0 ^~ inbuffer_data[712];
assign xnor1[713] = 1'b0 ^~ inbuffer_data[713];
assign xnor1[714] = 1'b0 ^~ inbuffer_data[714];
assign xnor1[715] = 1'b0 ^~ inbuffer_data[715];
assign xnor1[716] = 1'b0 ^~ inbuffer_data[716];
assign xnor1[717] = 1'b1 ^~ inbuffer_data[717];
assign xnor1[718] = 1'b0 ^~ inbuffer_data[718];
assign xnor1[719] = 1'b0 ^~ inbuffer_data[719];
assign xnor1[720] = 1'b1 ^~ inbuffer_data[720];
assign xnor1[721] = 1'b1 ^~ inbuffer_data[721];
assign xnor1[722] = 1'b1 ^~ inbuffer_data[722];
assign xnor1[723] = 1'b0 ^~ inbuffer_data[723];
assign xnor1[724] = 1'b1 ^~ inbuffer_data[724];
assign xnor1[725] = 1'b1 ^~ inbuffer_data[725];
assign xnor1[726] = 1'b0 ^~ inbuffer_data[726];
assign xnor1[727] = 1'b1 ^~ inbuffer_data[727];
assign xnor1[728] = 1'b1 ^~ inbuffer_data[728];
assign xnor1[729] = 1'b1 ^~ inbuffer_data[729];
assign xnor1[730] = 1'b0 ^~ inbuffer_data[730];
assign xnor1[731] = 1'b1 ^~ inbuffer_data[731];
assign xnor1[732] = 1'b0 ^~ inbuffer_data[732];
assign xnor1[733] = 1'b1 ^~ inbuffer_data[733];
assign xnor1[734] = 1'b1 ^~ inbuffer_data[734];
assign xnor1[735] = 1'b1 ^~ inbuffer_data[735];
assign xnor1[736] = 1'b0 ^~ inbuffer_data[736];
assign xnor1[737] = 1'b1 ^~ inbuffer_data[737];
assign xnor1[738] = 1'b1 ^~ inbuffer_data[738];
assign xnor1[739] = 1'b0 ^~ inbuffer_data[739];
assign xnor1[740] = 1'b0 ^~ inbuffer_data[740];
assign xnor1[741] = 1'b0 ^~ inbuffer_data[741];
assign xnor1[742] = 1'b0 ^~ inbuffer_data[742];
assign xnor1[743] = 1'b0 ^~ inbuffer_data[743];
assign xnor1[744] = 1'b0 ^~ inbuffer_data[744];
assign xnor1[745] = 1'b1 ^~ inbuffer_data[745];
assign xnor1[746] = 1'b1 ^~ inbuffer_data[746];
assign xnor1[747] = 1'b0 ^~ inbuffer_data[747];
assign xnor1[748] = 1'b0 ^~ inbuffer_data[748];
assign xnor1[749] = 1'b1 ^~ inbuffer_data[749];
assign xnor1[750] = 1'b1 ^~ inbuffer_data[750];
assign xnor1[751] = 1'b1 ^~ inbuffer_data[751];
assign xnor1[752] = 1'b1 ^~ inbuffer_data[752];
assign xnor1[753] = 1'b0 ^~ inbuffer_data[753];
assign xnor1[754] = 1'b0 ^~ inbuffer_data[754];
assign xnor1[755] = 1'b0 ^~ inbuffer_data[755];
assign xnor1[756] = 1'b1 ^~ inbuffer_data[756];
assign xnor1[757] = 1'b0 ^~ inbuffer_data[757];
assign xnor1[758] = 1'b0 ^~ inbuffer_data[758];
assign xnor1[759] = 1'b0 ^~ inbuffer_data[759];
assign xnor1[760] = 1'b1 ^~ inbuffer_data[760];
assign xnor1[761] = 1'b1 ^~ inbuffer_data[761];
assign xnor1[762] = 1'b1 ^~ inbuffer_data[762];
assign xnor1[763] = 1'b1 ^~ inbuffer_data[763];
assign xnor1[764] = 1'b1 ^~ inbuffer_data[764];
assign xnor1[765] = 1'b1 ^~ inbuffer_data[765];
assign xnor1[766] = 1'b1 ^~ inbuffer_data[766];
assign xnor1[767] = 1'b1 ^~ inbuffer_data[767];
assign xnor1[768] = 1'b1 ^~ inbuffer_data[768];
assign xnor1[769] = 1'b1 ^~ inbuffer_data[769];
assign xnor1[770] = 1'b1 ^~ inbuffer_data[770];
assign xnor1[771] = 1'b1 ^~ inbuffer_data[771];
assign xnor1[772] = 1'b0 ^~ inbuffer_data[772];
assign xnor1[773] = 1'b0 ^~ inbuffer_data[773];
assign xnor1[774] = 1'b1 ^~ inbuffer_data[774];
assign xnor1[775] = 1'b1 ^~ inbuffer_data[775];
assign xnor1[776] = 1'b0 ^~ inbuffer_data[776];
assign xnor1[777] = 1'b0 ^~ inbuffer_data[777];
assign xnor1[778] = 1'b1 ^~ inbuffer_data[778];
assign xnor1[779] = 1'b1 ^~ inbuffer_data[779];
assign xnor1[780] = 1'b0 ^~ inbuffer_data[780];
assign xnor1[781] = 1'b1 ^~ inbuffer_data[781];
assign xnor1[782] = 1'b0 ^~ inbuffer_data[782];
assign xnor1[783] = 1'b1 ^~ inbuffer_data[783];
assign xnor2[0] = 1'b0 ^~ inbuffer_data[0];
assign xnor2[1] = 1'b0 ^~ inbuffer_data[1];
assign xnor2[2] = 1'b0 ^~ inbuffer_data[2];
assign xnor2[3] = 1'b1 ^~ inbuffer_data[3];
assign xnor2[4] = 1'b0 ^~ inbuffer_data[4];
assign xnor2[5] = 1'b1 ^~ inbuffer_data[5];
assign xnor2[6] = 1'b0 ^~ inbuffer_data[6];
assign xnor2[7] = 1'b1 ^~ inbuffer_data[7];
assign xnor2[8] = 1'b0 ^~ inbuffer_data[8];
assign xnor2[9] = 1'b1 ^~ inbuffer_data[9];
assign xnor2[10] = 1'b0 ^~ inbuffer_data[10];
assign xnor2[11] = 1'b0 ^~ inbuffer_data[11];
assign xnor2[12] = 1'b1 ^~ inbuffer_data[12];
assign xnor2[13] = 1'b0 ^~ inbuffer_data[13];
assign xnor2[14] = 1'b0 ^~ inbuffer_data[14];
assign xnor2[15] = 1'b0 ^~ inbuffer_data[15];
assign xnor2[16] = 1'b0 ^~ inbuffer_data[16];
assign xnor2[17] = 1'b1 ^~ inbuffer_data[17];
assign xnor2[18] = 1'b0 ^~ inbuffer_data[18];
assign xnor2[19] = 1'b0 ^~ inbuffer_data[19];
assign xnor2[20] = 1'b0 ^~ inbuffer_data[20];
assign xnor2[21] = 1'b0 ^~ inbuffer_data[21];
assign xnor2[22] = 1'b1 ^~ inbuffer_data[22];
assign xnor2[23] = 1'b1 ^~ inbuffer_data[23];
assign xnor2[24] = 1'b1 ^~ inbuffer_data[24];
assign xnor2[25] = 1'b0 ^~ inbuffer_data[25];
assign xnor2[26] = 1'b1 ^~ inbuffer_data[26];
assign xnor2[27] = 1'b0 ^~ inbuffer_data[27];
assign xnor2[28] = 1'b1 ^~ inbuffer_data[28];
assign xnor2[29] = 1'b0 ^~ inbuffer_data[29];
assign xnor2[30] = 1'b0 ^~ inbuffer_data[30];
assign xnor2[31] = 1'b1 ^~ inbuffer_data[31];
assign xnor2[32] = 1'b0 ^~ inbuffer_data[32];
assign xnor2[33] = 1'b1 ^~ inbuffer_data[33];
assign xnor2[34] = 1'b0 ^~ inbuffer_data[34];
assign xnor2[35] = 1'b1 ^~ inbuffer_data[35];
assign xnor2[36] = 1'b1 ^~ inbuffer_data[36];
assign xnor2[37] = 1'b0 ^~ inbuffer_data[37];
assign xnor2[38] = 1'b0 ^~ inbuffer_data[38];
assign xnor2[39] = 1'b0 ^~ inbuffer_data[39];
assign xnor2[40] = 1'b0 ^~ inbuffer_data[40];
assign xnor2[41] = 1'b1 ^~ inbuffer_data[41];
assign xnor2[42] = 1'b0 ^~ inbuffer_data[42];
assign xnor2[43] = 1'b1 ^~ inbuffer_data[43];
assign xnor2[44] = 1'b1 ^~ inbuffer_data[44];
assign xnor2[45] = 1'b1 ^~ inbuffer_data[45];
assign xnor2[46] = 1'b1 ^~ inbuffer_data[46];
assign xnor2[47] = 1'b0 ^~ inbuffer_data[47];
assign xnor2[48] = 1'b1 ^~ inbuffer_data[48];
assign xnor2[49] = 1'b1 ^~ inbuffer_data[49];
assign xnor2[50] = 1'b0 ^~ inbuffer_data[50];
assign xnor2[51] = 1'b0 ^~ inbuffer_data[51];
assign xnor2[52] = 1'b0 ^~ inbuffer_data[52];
assign xnor2[53] = 1'b1 ^~ inbuffer_data[53];
assign xnor2[54] = 1'b0 ^~ inbuffer_data[54];
assign xnor2[55] = 1'b1 ^~ inbuffer_data[55];
assign xnor2[56] = 1'b0 ^~ inbuffer_data[56];
assign xnor2[57] = 1'b0 ^~ inbuffer_data[57];
assign xnor2[58] = 1'b0 ^~ inbuffer_data[58];
assign xnor2[59] = 1'b1 ^~ inbuffer_data[59];
assign xnor2[60] = 1'b0 ^~ inbuffer_data[60];
assign xnor2[61] = 1'b1 ^~ inbuffer_data[61];
assign xnor2[62] = 1'b1 ^~ inbuffer_data[62];
assign xnor2[63] = 1'b0 ^~ inbuffer_data[63];
assign xnor2[64] = 1'b1 ^~ inbuffer_data[64];
assign xnor2[65] = 1'b1 ^~ inbuffer_data[65];
assign xnor2[66] = 1'b1 ^~ inbuffer_data[66];
assign xnor2[67] = 1'b0 ^~ inbuffer_data[67];
assign xnor2[68] = 1'b1 ^~ inbuffer_data[68];
assign xnor2[69] = 1'b1 ^~ inbuffer_data[69];
assign xnor2[70] = 1'b1 ^~ inbuffer_data[70];
assign xnor2[71] = 1'b1 ^~ inbuffer_data[71];
assign xnor2[72] = 1'b0 ^~ inbuffer_data[72];
assign xnor2[73] = 1'b0 ^~ inbuffer_data[73];
assign xnor2[74] = 1'b0 ^~ inbuffer_data[74];
assign xnor2[75] = 1'b0 ^~ inbuffer_data[75];
assign xnor2[76] = 1'b1 ^~ inbuffer_data[76];
assign xnor2[77] = 1'b1 ^~ inbuffer_data[77];
assign xnor2[78] = 1'b1 ^~ inbuffer_data[78];
assign xnor2[79] = 1'b1 ^~ inbuffer_data[79];
assign xnor2[80] = 1'b0 ^~ inbuffer_data[80];
assign xnor2[81] = 1'b0 ^~ inbuffer_data[81];
assign xnor2[82] = 1'b1 ^~ inbuffer_data[82];
assign xnor2[83] = 1'b1 ^~ inbuffer_data[83];
assign xnor2[84] = 1'b0 ^~ inbuffer_data[84];
assign xnor2[85] = 1'b0 ^~ inbuffer_data[85];
assign xnor2[86] = 1'b0 ^~ inbuffer_data[86];
assign xnor2[87] = 1'b0 ^~ inbuffer_data[87];
assign xnor2[88] = 1'b0 ^~ inbuffer_data[88];
assign xnor2[89] = 1'b1 ^~ inbuffer_data[89];
assign xnor2[90] = 1'b1 ^~ inbuffer_data[90];
assign xnor2[91] = 1'b0 ^~ inbuffer_data[91];
assign xnor2[92] = 1'b0 ^~ inbuffer_data[92];
assign xnor2[93] = 1'b1 ^~ inbuffer_data[93];
assign xnor2[94] = 1'b1 ^~ inbuffer_data[94];
assign xnor2[95] = 1'b1 ^~ inbuffer_data[95];
assign xnor2[96] = 1'b1 ^~ inbuffer_data[96];
assign xnor2[97] = 1'b1 ^~ inbuffer_data[97];
assign xnor2[98] = 1'b1 ^~ inbuffer_data[98];
assign xnor2[99] = 1'b1 ^~ inbuffer_data[99];
assign xnor2[100] = 1'b1 ^~ inbuffer_data[100];
assign xnor2[101] = 1'b1 ^~ inbuffer_data[101];
assign xnor2[102] = 1'b0 ^~ inbuffer_data[102];
assign xnor2[103] = 1'b0 ^~ inbuffer_data[103];
assign xnor2[104] = 1'b0 ^~ inbuffer_data[104];
assign xnor2[105] = 1'b0 ^~ inbuffer_data[105];
assign xnor2[106] = 1'b0 ^~ inbuffer_data[106];
assign xnor2[107] = 1'b0 ^~ inbuffer_data[107];
assign xnor2[108] = 1'b0 ^~ inbuffer_data[108];
assign xnor2[109] = 1'b0 ^~ inbuffer_data[109];
assign xnor2[110] = 1'b1 ^~ inbuffer_data[110];
assign xnor2[111] = 1'b0 ^~ inbuffer_data[111];
assign xnor2[112] = 1'b1 ^~ inbuffer_data[112];
assign xnor2[113] = 1'b1 ^~ inbuffer_data[113];
assign xnor2[114] = 1'b0 ^~ inbuffer_data[114];
assign xnor2[115] = 1'b0 ^~ inbuffer_data[115];
assign xnor2[116] = 1'b0 ^~ inbuffer_data[116];
assign xnor2[117] = 1'b0 ^~ inbuffer_data[117];
assign xnor2[118] = 1'b1 ^~ inbuffer_data[118];
assign xnor2[119] = 1'b1 ^~ inbuffer_data[119];
assign xnor2[120] = 1'b1 ^~ inbuffer_data[120];
assign xnor2[121] = 1'b1 ^~ inbuffer_data[121];
assign xnor2[122] = 1'b1 ^~ inbuffer_data[122];
assign xnor2[123] = 1'b0 ^~ inbuffer_data[123];
assign xnor2[124] = 1'b1 ^~ inbuffer_data[124];
assign xnor2[125] = 1'b1 ^~ inbuffer_data[125];
assign xnor2[126] = 1'b1 ^~ inbuffer_data[126];
assign xnor2[127] = 1'b1 ^~ inbuffer_data[127];
assign xnor2[128] = 1'b1 ^~ inbuffer_data[128];
assign xnor2[129] = 1'b1 ^~ inbuffer_data[129];
assign xnor2[130] = 1'b1 ^~ inbuffer_data[130];
assign xnor2[131] = 1'b0 ^~ inbuffer_data[131];
assign xnor2[132] = 1'b0 ^~ inbuffer_data[132];
assign xnor2[133] = 1'b0 ^~ inbuffer_data[133];
assign xnor2[134] = 1'b0 ^~ inbuffer_data[134];
assign xnor2[135] = 1'b0 ^~ inbuffer_data[135];
assign xnor2[136] = 1'b0 ^~ inbuffer_data[136];
assign xnor2[137] = 1'b0 ^~ inbuffer_data[137];
assign xnor2[138] = 1'b0 ^~ inbuffer_data[138];
assign xnor2[139] = 1'b0 ^~ inbuffer_data[139];
assign xnor2[140] = 1'b0 ^~ inbuffer_data[140];
assign xnor2[141] = 1'b0 ^~ inbuffer_data[141];
assign xnor2[142] = 1'b0 ^~ inbuffer_data[142];
assign xnor2[143] = 1'b0 ^~ inbuffer_data[143];
assign xnor2[144] = 1'b0 ^~ inbuffer_data[144];
assign xnor2[145] = 1'b0 ^~ inbuffer_data[145];
assign xnor2[146] = 1'b1 ^~ inbuffer_data[146];
assign xnor2[147] = 1'b1 ^~ inbuffer_data[147];
assign xnor2[148] = 1'b1 ^~ inbuffer_data[148];
assign xnor2[149] = 1'b1 ^~ inbuffer_data[149];
assign xnor2[150] = 1'b1 ^~ inbuffer_data[150];
assign xnor2[151] = 1'b1 ^~ inbuffer_data[151];
assign xnor2[152] = 1'b1 ^~ inbuffer_data[152];
assign xnor2[153] = 1'b1 ^~ inbuffer_data[153];
assign xnor2[154] = 1'b1 ^~ inbuffer_data[154];
assign xnor2[155] = 1'b1 ^~ inbuffer_data[155];
assign xnor2[156] = 1'b1 ^~ inbuffer_data[156];
assign xnor2[157] = 1'b1 ^~ inbuffer_data[157];
assign xnor2[158] = 1'b1 ^~ inbuffer_data[158];
assign xnor2[159] = 1'b0 ^~ inbuffer_data[159];
assign xnor2[160] = 1'b1 ^~ inbuffer_data[160];
assign xnor2[161] = 1'b0 ^~ inbuffer_data[161];
assign xnor2[162] = 1'b1 ^~ inbuffer_data[162];
assign xnor2[163] = 1'b0 ^~ inbuffer_data[163];
assign xnor2[164] = 1'b0 ^~ inbuffer_data[164];
assign xnor2[165] = 1'b0 ^~ inbuffer_data[165];
assign xnor2[166] = 1'b1 ^~ inbuffer_data[166];
assign xnor2[167] = 1'b1 ^~ inbuffer_data[167];
assign xnor2[168] = 1'b1 ^~ inbuffer_data[168];
assign xnor2[169] = 1'b0 ^~ inbuffer_data[169];
assign xnor2[170] = 1'b1 ^~ inbuffer_data[170];
assign xnor2[171] = 1'b1 ^~ inbuffer_data[171];
assign xnor2[172] = 1'b0 ^~ inbuffer_data[172];
assign xnor2[173] = 1'b1 ^~ inbuffer_data[173];
assign xnor2[174] = 1'b1 ^~ inbuffer_data[174];
assign xnor2[175] = 1'b1 ^~ inbuffer_data[175];
assign xnor2[176] = 1'b1 ^~ inbuffer_data[176];
assign xnor2[177] = 1'b1 ^~ inbuffer_data[177];
assign xnor2[178] = 1'b1 ^~ inbuffer_data[178];
assign xnor2[179] = 1'b1 ^~ inbuffer_data[179];
assign xnor2[180] = 1'b1 ^~ inbuffer_data[180];
assign xnor2[181] = 1'b1 ^~ inbuffer_data[181];
assign xnor2[182] = 1'b1 ^~ inbuffer_data[182];
assign xnor2[183] = 1'b1 ^~ inbuffer_data[183];
assign xnor2[184] = 1'b1 ^~ inbuffer_data[184];
assign xnor2[185] = 1'b0 ^~ inbuffer_data[185];
assign xnor2[186] = 1'b1 ^~ inbuffer_data[186];
assign xnor2[187] = 1'b1 ^~ inbuffer_data[187];
assign xnor2[188] = 1'b0 ^~ inbuffer_data[188];
assign xnor2[189] = 1'b0 ^~ inbuffer_data[189];
assign xnor2[190] = 1'b0 ^~ inbuffer_data[190];
assign xnor2[191] = 1'b0 ^~ inbuffer_data[191];
assign xnor2[192] = 1'b0 ^~ inbuffer_data[192];
assign xnor2[193] = 1'b1 ^~ inbuffer_data[193];
assign xnor2[194] = 1'b1 ^~ inbuffer_data[194];
assign xnor2[195] = 1'b0 ^~ inbuffer_data[195];
assign xnor2[196] = 1'b0 ^~ inbuffer_data[196];
assign xnor2[197] = 1'b0 ^~ inbuffer_data[197];
assign xnor2[198] = 1'b0 ^~ inbuffer_data[198];
assign xnor2[199] = 1'b1 ^~ inbuffer_data[199];
assign xnor2[200] = 1'b1 ^~ inbuffer_data[200];
assign xnor2[201] = 1'b1 ^~ inbuffer_data[201];
assign xnor2[202] = 1'b1 ^~ inbuffer_data[202];
assign xnor2[203] = 1'b0 ^~ inbuffer_data[203];
assign xnor2[204] = 1'b1 ^~ inbuffer_data[204];
assign xnor2[205] = 1'b1 ^~ inbuffer_data[205];
assign xnor2[206] = 1'b1 ^~ inbuffer_data[206];
assign xnor2[207] = 1'b1 ^~ inbuffer_data[207];
assign xnor2[208] = 1'b1 ^~ inbuffer_data[208];
assign xnor2[209] = 1'b0 ^~ inbuffer_data[209];
assign xnor2[210] = 1'b1 ^~ inbuffer_data[210];
assign xnor2[211] = 1'b1 ^~ inbuffer_data[211];
assign xnor2[212] = 1'b1 ^~ inbuffer_data[212];
assign xnor2[213] = 1'b0 ^~ inbuffer_data[213];
assign xnor2[214] = 1'b0 ^~ inbuffer_data[214];
assign xnor2[215] = 1'b1 ^~ inbuffer_data[215];
assign xnor2[216] = 1'b0 ^~ inbuffer_data[216];
assign xnor2[217] = 1'b1 ^~ inbuffer_data[217];
assign xnor2[218] = 1'b1 ^~ inbuffer_data[218];
assign xnor2[219] = 1'b0 ^~ inbuffer_data[219];
assign xnor2[220] = 1'b0 ^~ inbuffer_data[220];
assign xnor2[221] = 1'b0 ^~ inbuffer_data[221];
assign xnor2[222] = 1'b1 ^~ inbuffer_data[222];
assign xnor2[223] = 1'b1 ^~ inbuffer_data[223];
assign xnor2[224] = 1'b0 ^~ inbuffer_data[224];
assign xnor2[225] = 1'b0 ^~ inbuffer_data[225];
assign xnor2[226] = 1'b1 ^~ inbuffer_data[226];
assign xnor2[227] = 1'b1 ^~ inbuffer_data[227];
assign xnor2[228] = 1'b1 ^~ inbuffer_data[228];
assign xnor2[229] = 1'b0 ^~ inbuffer_data[229];
assign xnor2[230] = 1'b1 ^~ inbuffer_data[230];
assign xnor2[231] = 1'b1 ^~ inbuffer_data[231];
assign xnor2[232] = 1'b1 ^~ inbuffer_data[232];
assign xnor2[233] = 1'b0 ^~ inbuffer_data[233];
assign xnor2[234] = 1'b1 ^~ inbuffer_data[234];
assign xnor2[235] = 1'b1 ^~ inbuffer_data[235];
assign xnor2[236] = 1'b0 ^~ inbuffer_data[236];
assign xnor2[237] = 1'b0 ^~ inbuffer_data[237];
assign xnor2[238] = 1'b1 ^~ inbuffer_data[238];
assign xnor2[239] = 1'b1 ^~ inbuffer_data[239];
assign xnor2[240] = 1'b1 ^~ inbuffer_data[240];
assign xnor2[241] = 1'b1 ^~ inbuffer_data[241];
assign xnor2[242] = 1'b0 ^~ inbuffer_data[242];
assign xnor2[243] = 1'b1 ^~ inbuffer_data[243];
assign xnor2[244] = 1'b1 ^~ inbuffer_data[244];
assign xnor2[245] = 1'b0 ^~ inbuffer_data[245];
assign xnor2[246] = 1'b1 ^~ inbuffer_data[246];
assign xnor2[247] = 1'b0 ^~ inbuffer_data[247];
assign xnor2[248] = 1'b0 ^~ inbuffer_data[248];
assign xnor2[249] = 1'b0 ^~ inbuffer_data[249];
assign xnor2[250] = 1'b0 ^~ inbuffer_data[250];
assign xnor2[251] = 1'b0 ^~ inbuffer_data[251];
assign xnor2[252] = 1'b1 ^~ inbuffer_data[252];
assign xnor2[253] = 1'b1 ^~ inbuffer_data[253];
assign xnor2[254] = 1'b1 ^~ inbuffer_data[254];
assign xnor2[255] = 1'b0 ^~ inbuffer_data[255];
assign xnor2[256] = 1'b1 ^~ inbuffer_data[256];
assign xnor2[257] = 1'b1 ^~ inbuffer_data[257];
assign xnor2[258] = 1'b0 ^~ inbuffer_data[258];
assign xnor2[259] = 1'b0 ^~ inbuffer_data[259];
assign xnor2[260] = 1'b1 ^~ inbuffer_data[260];
assign xnor2[261] = 1'b1 ^~ inbuffer_data[261];
assign xnor2[262] = 1'b0 ^~ inbuffer_data[262];
assign xnor2[263] = 1'b1 ^~ inbuffer_data[263];
assign xnor2[264] = 1'b1 ^~ inbuffer_data[264];
assign xnor2[265] = 1'b0 ^~ inbuffer_data[265];
assign xnor2[266] = 1'b1 ^~ inbuffer_data[266];
assign xnor2[267] = 1'b1 ^~ inbuffer_data[267];
assign xnor2[268] = 1'b1 ^~ inbuffer_data[268];
assign xnor2[269] = 1'b1 ^~ inbuffer_data[269];
assign xnor2[270] = 1'b1 ^~ inbuffer_data[270];
assign xnor2[271] = 1'b1 ^~ inbuffer_data[271];
assign xnor2[272] = 1'b0 ^~ inbuffer_data[272];
assign xnor2[273] = 1'b0 ^~ inbuffer_data[273];
assign xnor2[274] = 1'b1 ^~ inbuffer_data[274];
assign xnor2[275] = 1'b0 ^~ inbuffer_data[275];
assign xnor2[276] = 1'b0 ^~ inbuffer_data[276];
assign xnor2[277] = 1'b0 ^~ inbuffer_data[277];
assign xnor2[278] = 1'b0 ^~ inbuffer_data[278];
assign xnor2[279] = 1'b1 ^~ inbuffer_data[279];
assign xnor2[280] = 1'b1 ^~ inbuffer_data[280];
assign xnor2[281] = 1'b0 ^~ inbuffer_data[281];
assign xnor2[282] = 1'b0 ^~ inbuffer_data[282];
assign xnor2[283] = 1'b0 ^~ inbuffer_data[283];
assign xnor2[284] = 1'b0 ^~ inbuffer_data[284];
assign xnor2[285] = 1'b1 ^~ inbuffer_data[285];
assign xnor2[286] = 1'b1 ^~ inbuffer_data[286];
assign xnor2[287] = 1'b0 ^~ inbuffer_data[287];
assign xnor2[288] = 1'b0 ^~ inbuffer_data[288];
assign xnor2[289] = 1'b0 ^~ inbuffer_data[289];
assign xnor2[290] = 1'b0 ^~ inbuffer_data[290];
assign xnor2[291] = 1'b0 ^~ inbuffer_data[291];
assign xnor2[292] = 1'b0 ^~ inbuffer_data[292];
assign xnor2[293] = 1'b0 ^~ inbuffer_data[293];
assign xnor2[294] = 1'b0 ^~ inbuffer_data[294];
assign xnor2[295] = 1'b0 ^~ inbuffer_data[295];
assign xnor2[296] = 1'b0 ^~ inbuffer_data[296];
assign xnor2[297] = 1'b1 ^~ inbuffer_data[297];
assign xnor2[298] = 1'b1 ^~ inbuffer_data[298];
assign xnor2[299] = 1'b0 ^~ inbuffer_data[299];
assign xnor2[300] = 1'b1 ^~ inbuffer_data[300];
assign xnor2[301] = 1'b1 ^~ inbuffer_data[301];
assign xnor2[302] = 1'b0 ^~ inbuffer_data[302];
assign xnor2[303] = 1'b0 ^~ inbuffer_data[303];
assign xnor2[304] = 1'b0 ^~ inbuffer_data[304];
assign xnor2[305] = 1'b0 ^~ inbuffer_data[305];
assign xnor2[306] = 1'b1 ^~ inbuffer_data[306];
assign xnor2[307] = 1'b0 ^~ inbuffer_data[307];
assign xnor2[308] = 1'b0 ^~ inbuffer_data[308];
assign xnor2[309] = 1'b0 ^~ inbuffer_data[309];
assign xnor2[310] = 1'b1 ^~ inbuffer_data[310];
assign xnor2[311] = 1'b0 ^~ inbuffer_data[311];
assign xnor2[312] = 1'b1 ^~ inbuffer_data[312];
assign xnor2[313] = 1'b0 ^~ inbuffer_data[313];
assign xnor2[314] = 1'b0 ^~ inbuffer_data[314];
assign xnor2[315] = 1'b0 ^~ inbuffer_data[315];
assign xnor2[316] = 1'b0 ^~ inbuffer_data[316];
assign xnor2[317] = 1'b0 ^~ inbuffer_data[317];
assign xnor2[318] = 1'b0 ^~ inbuffer_data[318];
assign xnor2[319] = 1'b0 ^~ inbuffer_data[319];
assign xnor2[320] = 1'b0 ^~ inbuffer_data[320];
assign xnor2[321] = 1'b0 ^~ inbuffer_data[321];
assign xnor2[322] = 1'b0 ^~ inbuffer_data[322];
assign xnor2[323] = 1'b0 ^~ inbuffer_data[323];
assign xnor2[324] = 1'b0 ^~ inbuffer_data[324];
assign xnor2[325] = 1'b0 ^~ inbuffer_data[325];
assign xnor2[326] = 1'b0 ^~ inbuffer_data[326];
assign xnor2[327] = 1'b1 ^~ inbuffer_data[327];
assign xnor2[328] = 1'b1 ^~ inbuffer_data[328];
assign xnor2[329] = 1'b0 ^~ inbuffer_data[329];
assign xnor2[330] = 1'b1 ^~ inbuffer_data[330];
assign xnor2[331] = 1'b0 ^~ inbuffer_data[331];
assign xnor2[332] = 1'b0 ^~ inbuffer_data[332];
assign xnor2[333] = 1'b1 ^~ inbuffer_data[333];
assign xnor2[334] = 1'b0 ^~ inbuffer_data[334];
assign xnor2[335] = 1'b1 ^~ inbuffer_data[335];
assign xnor2[336] = 1'b0 ^~ inbuffer_data[336];
assign xnor2[337] = 1'b0 ^~ inbuffer_data[337];
assign xnor2[338] = 1'b1 ^~ inbuffer_data[338];
assign xnor2[339] = 1'b1 ^~ inbuffer_data[339];
assign xnor2[340] = 1'b0 ^~ inbuffer_data[340];
assign xnor2[341] = 1'b0 ^~ inbuffer_data[341];
assign xnor2[342] = 1'b0 ^~ inbuffer_data[342];
assign xnor2[343] = 1'b0 ^~ inbuffer_data[343];
assign xnor2[344] = 1'b0 ^~ inbuffer_data[344];
assign xnor2[345] = 1'b0 ^~ inbuffer_data[345];
assign xnor2[346] = 1'b0 ^~ inbuffer_data[346];
assign xnor2[347] = 1'b0 ^~ inbuffer_data[347];
assign xnor2[348] = 1'b0 ^~ inbuffer_data[348];
assign xnor2[349] = 1'b0 ^~ inbuffer_data[349];
assign xnor2[350] = 1'b0 ^~ inbuffer_data[350];
assign xnor2[351] = 1'b0 ^~ inbuffer_data[351];
assign xnor2[352] = 1'b0 ^~ inbuffer_data[352];
assign xnor2[353] = 1'b0 ^~ inbuffer_data[353];
assign xnor2[354] = 1'b0 ^~ inbuffer_data[354];
assign xnor2[355] = 1'b1 ^~ inbuffer_data[355];
assign xnor2[356] = 1'b1 ^~ inbuffer_data[356];
assign xnor2[357] = 1'b1 ^~ inbuffer_data[357];
assign xnor2[358] = 1'b0 ^~ inbuffer_data[358];
assign xnor2[359] = 1'b0 ^~ inbuffer_data[359];
assign xnor2[360] = 1'b0 ^~ inbuffer_data[360];
assign xnor2[361] = 1'b1 ^~ inbuffer_data[361];
assign xnor2[362] = 1'b1 ^~ inbuffer_data[362];
assign xnor2[363] = 1'b1 ^~ inbuffer_data[363];
assign xnor2[364] = 1'b1 ^~ inbuffer_data[364];
assign xnor2[365] = 1'b0 ^~ inbuffer_data[365];
assign xnor2[366] = 1'b0 ^~ inbuffer_data[366];
assign xnor2[367] = 1'b0 ^~ inbuffer_data[367];
assign xnor2[368] = 1'b0 ^~ inbuffer_data[368];
assign xnor2[369] = 1'b0 ^~ inbuffer_data[369];
assign xnor2[370] = 1'b0 ^~ inbuffer_data[370];
assign xnor2[371] = 1'b0 ^~ inbuffer_data[371];
assign xnor2[372] = 1'b0 ^~ inbuffer_data[372];
assign xnor2[373] = 1'b0 ^~ inbuffer_data[373];
assign xnor2[374] = 1'b0 ^~ inbuffer_data[374];
assign xnor2[375] = 1'b0 ^~ inbuffer_data[375];
assign xnor2[376] = 1'b0 ^~ inbuffer_data[376];
assign xnor2[377] = 1'b0 ^~ inbuffer_data[377];
assign xnor2[378] = 1'b0 ^~ inbuffer_data[378];
assign xnor2[379] = 1'b0 ^~ inbuffer_data[379];
assign xnor2[380] = 1'b1 ^~ inbuffer_data[380];
assign xnor2[381] = 1'b0 ^~ inbuffer_data[381];
assign xnor2[382] = 1'b0 ^~ inbuffer_data[382];
assign xnor2[383] = 1'b0 ^~ inbuffer_data[383];
assign xnor2[384] = 1'b0 ^~ inbuffer_data[384];
assign xnor2[385] = 1'b0 ^~ inbuffer_data[385];
assign xnor2[386] = 1'b0 ^~ inbuffer_data[386];
assign xnor2[387] = 1'b0 ^~ inbuffer_data[387];
assign xnor2[388] = 1'b1 ^~ inbuffer_data[388];
assign xnor2[389] = 1'b1 ^~ inbuffer_data[389];
assign xnor2[390] = 1'b1 ^~ inbuffer_data[390];
assign xnor2[391] = 1'b1 ^~ inbuffer_data[391];
assign xnor2[392] = 1'b1 ^~ inbuffer_data[392];
assign xnor2[393] = 1'b1 ^~ inbuffer_data[393];
assign xnor2[394] = 1'b0 ^~ inbuffer_data[394];
assign xnor2[395] = 1'b0 ^~ inbuffer_data[395];
assign xnor2[396] = 1'b0 ^~ inbuffer_data[396];
assign xnor2[397] = 1'b0 ^~ inbuffer_data[397];
assign xnor2[398] = 1'b0 ^~ inbuffer_data[398];
assign xnor2[399] = 1'b0 ^~ inbuffer_data[399];
assign xnor2[400] = 1'b0 ^~ inbuffer_data[400];
assign xnor2[401] = 1'b0 ^~ inbuffer_data[401];
assign xnor2[402] = 1'b0 ^~ inbuffer_data[402];
assign xnor2[403] = 1'b0 ^~ inbuffer_data[403];
assign xnor2[404] = 1'b1 ^~ inbuffer_data[404];
assign xnor2[405] = 1'b1 ^~ inbuffer_data[405];
assign xnor2[406] = 1'b1 ^~ inbuffer_data[406];
assign xnor2[407] = 1'b1 ^~ inbuffer_data[407];
assign xnor2[408] = 1'b1 ^~ inbuffer_data[408];
assign xnor2[409] = 1'b0 ^~ inbuffer_data[409];
assign xnor2[410] = 1'b0 ^~ inbuffer_data[410];
assign xnor2[411] = 1'b0 ^~ inbuffer_data[411];
assign xnor2[412] = 1'b1 ^~ inbuffer_data[412];
assign xnor2[413] = 1'b0 ^~ inbuffer_data[413];
assign xnor2[414] = 1'b0 ^~ inbuffer_data[414];
assign xnor2[415] = 1'b1 ^~ inbuffer_data[415];
assign xnor2[416] = 1'b0 ^~ inbuffer_data[416];
assign xnor2[417] = 1'b1 ^~ inbuffer_data[417];
assign xnor2[418] = 1'b1 ^~ inbuffer_data[418];
assign xnor2[419] = 1'b0 ^~ inbuffer_data[419];
assign xnor2[420] = 1'b1 ^~ inbuffer_data[420];
assign xnor2[421] = 1'b0 ^~ inbuffer_data[421];
assign xnor2[422] = 1'b0 ^~ inbuffer_data[422];
assign xnor2[423] = 1'b0 ^~ inbuffer_data[423];
assign xnor2[424] = 1'b1 ^~ inbuffer_data[424];
assign xnor2[425] = 1'b0 ^~ inbuffer_data[425];
assign xnor2[426] = 1'b1 ^~ inbuffer_data[426];
assign xnor2[427] = 1'b0 ^~ inbuffer_data[427];
assign xnor2[428] = 1'b1 ^~ inbuffer_data[428];
assign xnor2[429] = 1'b1 ^~ inbuffer_data[429];
assign xnor2[430] = 1'b1 ^~ inbuffer_data[430];
assign xnor2[431] = 1'b0 ^~ inbuffer_data[431];
assign xnor2[432] = 1'b1 ^~ inbuffer_data[432];
assign xnor2[433] = 1'b1 ^~ inbuffer_data[433];
assign xnor2[434] = 1'b0 ^~ inbuffer_data[434];
assign xnor2[435] = 1'b1 ^~ inbuffer_data[435];
assign xnor2[436] = 1'b1 ^~ inbuffer_data[436];
assign xnor2[437] = 1'b0 ^~ inbuffer_data[437];
assign xnor2[438] = 1'b0 ^~ inbuffer_data[438];
assign xnor2[439] = 1'b1 ^~ inbuffer_data[439];
assign xnor2[440] = 1'b0 ^~ inbuffer_data[440];
assign xnor2[441] = 1'b0 ^~ inbuffer_data[441];
assign xnor2[442] = 1'b0 ^~ inbuffer_data[442];
assign xnor2[443] = 1'b0 ^~ inbuffer_data[443];
assign xnor2[444] = 1'b1 ^~ inbuffer_data[444];
assign xnor2[445] = 1'b1 ^~ inbuffer_data[445];
assign xnor2[446] = 1'b1 ^~ inbuffer_data[446];
assign xnor2[447] = 1'b1 ^~ inbuffer_data[447];
assign xnor2[448] = 1'b0 ^~ inbuffer_data[448];
assign xnor2[449] = 1'b0 ^~ inbuffer_data[449];
assign xnor2[450] = 1'b0 ^~ inbuffer_data[450];
assign xnor2[451] = 1'b1 ^~ inbuffer_data[451];
assign xnor2[452] = 1'b1 ^~ inbuffer_data[452];
assign xnor2[453] = 1'b1 ^~ inbuffer_data[453];
assign xnor2[454] = 1'b1 ^~ inbuffer_data[454];
assign xnor2[455] = 1'b1 ^~ inbuffer_data[455];
assign xnor2[456] = 1'b1 ^~ inbuffer_data[456];
assign xnor2[457] = 1'b1 ^~ inbuffer_data[457];
assign xnor2[458] = 1'b1 ^~ inbuffer_data[458];
assign xnor2[459] = 1'b1 ^~ inbuffer_data[459];
assign xnor2[460] = 1'b1 ^~ inbuffer_data[460];
assign xnor2[461] = 1'b1 ^~ inbuffer_data[461];
assign xnor2[462] = 1'b1 ^~ inbuffer_data[462];
assign xnor2[463] = 1'b1 ^~ inbuffer_data[463];
assign xnor2[464] = 1'b0 ^~ inbuffer_data[464];
assign xnor2[465] = 1'b1 ^~ inbuffer_data[465];
assign xnor2[466] = 1'b1 ^~ inbuffer_data[466];
assign xnor2[467] = 1'b0 ^~ inbuffer_data[467];
assign xnor2[468] = 1'b1 ^~ inbuffer_data[468];
assign xnor2[469] = 1'b1 ^~ inbuffer_data[469];
assign xnor2[470] = 1'b1 ^~ inbuffer_data[470];
assign xnor2[471] = 1'b1 ^~ inbuffer_data[471];
assign xnor2[472] = 1'b1 ^~ inbuffer_data[472];
assign xnor2[473] = 1'b1 ^~ inbuffer_data[473];
assign xnor2[474] = 1'b1 ^~ inbuffer_data[474];
assign xnor2[475] = 1'b0 ^~ inbuffer_data[475];
assign xnor2[476] = 1'b0 ^~ inbuffer_data[476];
assign xnor2[477] = 1'b1 ^~ inbuffer_data[477];
assign xnor2[478] = 1'b0 ^~ inbuffer_data[478];
assign xnor2[479] = 1'b1 ^~ inbuffer_data[479];
assign xnor2[480] = 1'b1 ^~ inbuffer_data[480];
assign xnor2[481] = 1'b1 ^~ inbuffer_data[481];
assign xnor2[482] = 1'b1 ^~ inbuffer_data[482];
assign xnor2[483] = 1'b1 ^~ inbuffer_data[483];
assign xnor2[484] = 1'b1 ^~ inbuffer_data[484];
assign xnor2[485] = 1'b1 ^~ inbuffer_data[485];
assign xnor2[486] = 1'b1 ^~ inbuffer_data[486];
assign xnor2[487] = 1'b1 ^~ inbuffer_data[487];
assign xnor2[488] = 1'b1 ^~ inbuffer_data[488];
assign xnor2[489] = 1'b1 ^~ inbuffer_data[489];
assign xnor2[490] = 1'b0 ^~ inbuffer_data[490];
assign xnor2[491] = 1'b1 ^~ inbuffer_data[491];
assign xnor2[492] = 1'b1 ^~ inbuffer_data[492];
assign xnor2[493] = 1'b0 ^~ inbuffer_data[493];
assign xnor2[494] = 1'b1 ^~ inbuffer_data[494];
assign xnor2[495] = 1'b0 ^~ inbuffer_data[495];
assign xnor2[496] = 1'b1 ^~ inbuffer_data[496];
assign xnor2[497] = 1'b0 ^~ inbuffer_data[497];
assign xnor2[498] = 1'b1 ^~ inbuffer_data[498];
assign xnor2[499] = 1'b1 ^~ inbuffer_data[499];
assign xnor2[500] = 1'b1 ^~ inbuffer_data[500];
assign xnor2[501] = 1'b1 ^~ inbuffer_data[501];
assign xnor2[502] = 1'b1 ^~ inbuffer_data[502];
assign xnor2[503] = 1'b0 ^~ inbuffer_data[503];
assign xnor2[504] = 1'b0 ^~ inbuffer_data[504];
assign xnor2[505] = 1'b1 ^~ inbuffer_data[505];
assign xnor2[506] = 1'b0 ^~ inbuffer_data[506];
assign xnor2[507] = 1'b1 ^~ inbuffer_data[507];
assign xnor2[508] = 1'b1 ^~ inbuffer_data[508];
assign xnor2[509] = 1'b1 ^~ inbuffer_data[509];
assign xnor2[510] = 1'b1 ^~ inbuffer_data[510];
assign xnor2[511] = 1'b1 ^~ inbuffer_data[511];
assign xnor2[512] = 1'b1 ^~ inbuffer_data[512];
assign xnor2[513] = 1'b1 ^~ inbuffer_data[513];
assign xnor2[514] = 1'b1 ^~ inbuffer_data[514];
assign xnor2[515] = 1'b1 ^~ inbuffer_data[515];
assign xnor2[516] = 1'b1 ^~ inbuffer_data[516];
assign xnor2[517] = 1'b1 ^~ inbuffer_data[517];
assign xnor2[518] = 1'b1 ^~ inbuffer_data[518];
assign xnor2[519] = 1'b0 ^~ inbuffer_data[519];
assign xnor2[520] = 1'b1 ^~ inbuffer_data[520];
assign xnor2[521] = 1'b1 ^~ inbuffer_data[521];
assign xnor2[522] = 1'b1 ^~ inbuffer_data[522];
assign xnor2[523] = 1'b1 ^~ inbuffer_data[523];
assign xnor2[524] = 1'b0 ^~ inbuffer_data[524];
assign xnor2[525] = 1'b0 ^~ inbuffer_data[525];
assign xnor2[526] = 1'b1 ^~ inbuffer_data[526];
assign xnor2[527] = 1'b1 ^~ inbuffer_data[527];
assign xnor2[528] = 1'b1 ^~ inbuffer_data[528];
assign xnor2[529] = 1'b1 ^~ inbuffer_data[529];
assign xnor2[530] = 1'b1 ^~ inbuffer_data[530];
assign xnor2[531] = 1'b1 ^~ inbuffer_data[531];
assign xnor2[532] = 1'b0 ^~ inbuffer_data[532];
assign xnor2[533] = 1'b0 ^~ inbuffer_data[533];
assign xnor2[534] = 1'b0 ^~ inbuffer_data[534];
assign xnor2[535] = 1'b0 ^~ inbuffer_data[535];
assign xnor2[536] = 1'b1 ^~ inbuffer_data[536];
assign xnor2[537] = 1'b1 ^~ inbuffer_data[537];
assign xnor2[538] = 1'b1 ^~ inbuffer_data[538];
assign xnor2[539] = 1'b1 ^~ inbuffer_data[539];
assign xnor2[540] = 1'b1 ^~ inbuffer_data[540];
assign xnor2[541] = 1'b1 ^~ inbuffer_data[541];
assign xnor2[542] = 1'b1 ^~ inbuffer_data[542];
assign xnor2[543] = 1'b1 ^~ inbuffer_data[543];
assign xnor2[544] = 1'b1 ^~ inbuffer_data[544];
assign xnor2[545] = 1'b1 ^~ inbuffer_data[545];
assign xnor2[546] = 1'b1 ^~ inbuffer_data[546];
assign xnor2[547] = 1'b1 ^~ inbuffer_data[547];
assign xnor2[548] = 1'b0 ^~ inbuffer_data[548];
assign xnor2[549] = 1'b1 ^~ inbuffer_data[549];
assign xnor2[550] = 1'b0 ^~ inbuffer_data[550];
assign xnor2[551] = 1'b1 ^~ inbuffer_data[551];
assign xnor2[552] = 1'b1 ^~ inbuffer_data[552];
assign xnor2[553] = 1'b1 ^~ inbuffer_data[553];
assign xnor2[554] = 1'b1 ^~ inbuffer_data[554];
assign xnor2[555] = 1'b1 ^~ inbuffer_data[555];
assign xnor2[556] = 1'b1 ^~ inbuffer_data[556];
assign xnor2[557] = 1'b1 ^~ inbuffer_data[557];
assign xnor2[558] = 1'b1 ^~ inbuffer_data[558];
assign xnor2[559] = 1'b1 ^~ inbuffer_data[559];
assign xnor2[560] = 1'b0 ^~ inbuffer_data[560];
assign xnor2[561] = 1'b1 ^~ inbuffer_data[561];
assign xnor2[562] = 1'b1 ^~ inbuffer_data[562];
assign xnor2[563] = 1'b0 ^~ inbuffer_data[563];
assign xnor2[564] = 1'b1 ^~ inbuffer_data[564];
assign xnor2[565] = 1'b1 ^~ inbuffer_data[565];
assign xnor2[566] = 1'b1 ^~ inbuffer_data[566];
assign xnor2[567] = 1'b1 ^~ inbuffer_data[567];
assign xnor2[568] = 1'b1 ^~ inbuffer_data[568];
assign xnor2[569] = 1'b1 ^~ inbuffer_data[569];
assign xnor2[570] = 1'b1 ^~ inbuffer_data[570];
assign xnor2[571] = 1'b1 ^~ inbuffer_data[571];
assign xnor2[572] = 1'b1 ^~ inbuffer_data[572];
assign xnor2[573] = 1'b0 ^~ inbuffer_data[573];
assign xnor2[574] = 1'b0 ^~ inbuffer_data[574];
assign xnor2[575] = 1'b1 ^~ inbuffer_data[575];
assign xnor2[576] = 1'b1 ^~ inbuffer_data[576];
assign xnor2[577] = 1'b0 ^~ inbuffer_data[577];
assign xnor2[578] = 1'b1 ^~ inbuffer_data[578];
assign xnor2[579] = 1'b1 ^~ inbuffer_data[579];
assign xnor2[580] = 1'b1 ^~ inbuffer_data[580];
assign xnor2[581] = 1'b1 ^~ inbuffer_data[581];
assign xnor2[582] = 1'b1 ^~ inbuffer_data[582];
assign xnor2[583] = 1'b1 ^~ inbuffer_data[583];
assign xnor2[584] = 1'b1 ^~ inbuffer_data[584];
assign xnor2[585] = 1'b0 ^~ inbuffer_data[585];
assign xnor2[586] = 1'b1 ^~ inbuffer_data[586];
assign xnor2[587] = 1'b0 ^~ inbuffer_data[587];
assign xnor2[588] = 1'b0 ^~ inbuffer_data[588];
assign xnor2[589] = 1'b0 ^~ inbuffer_data[589];
assign xnor2[590] = 1'b0 ^~ inbuffer_data[590];
assign xnor2[591] = 1'b1 ^~ inbuffer_data[591];
assign xnor2[592] = 1'b1 ^~ inbuffer_data[592];
assign xnor2[593] = 1'b1 ^~ inbuffer_data[593];
assign xnor2[594] = 1'b1 ^~ inbuffer_data[594];
assign xnor2[595] = 1'b1 ^~ inbuffer_data[595];
assign xnor2[596] = 1'b1 ^~ inbuffer_data[596];
assign xnor2[597] = 1'b1 ^~ inbuffer_data[597];
assign xnor2[598] = 1'b1 ^~ inbuffer_data[598];
assign xnor2[599] = 1'b1 ^~ inbuffer_data[599];
assign xnor2[600] = 1'b1 ^~ inbuffer_data[600];
assign xnor2[601] = 1'b0 ^~ inbuffer_data[601];
assign xnor2[602] = 1'b0 ^~ inbuffer_data[602];
assign xnor2[603] = 1'b0 ^~ inbuffer_data[603];
assign xnor2[604] = 1'b1 ^~ inbuffer_data[604];
assign xnor2[605] = 1'b1 ^~ inbuffer_data[605];
assign xnor2[606] = 1'b1 ^~ inbuffer_data[606];
assign xnor2[607] = 1'b1 ^~ inbuffer_data[607];
assign xnor2[608] = 1'b1 ^~ inbuffer_data[608];
assign xnor2[609] = 1'b1 ^~ inbuffer_data[609];
assign xnor2[610] = 1'b1 ^~ inbuffer_data[610];
assign xnor2[611] = 1'b1 ^~ inbuffer_data[611];
assign xnor2[612] = 1'b1 ^~ inbuffer_data[612];
assign xnor2[613] = 1'b1 ^~ inbuffer_data[613];
assign xnor2[614] = 1'b0 ^~ inbuffer_data[614];
assign xnor2[615] = 1'b0 ^~ inbuffer_data[615];
assign xnor2[616] = 1'b1 ^~ inbuffer_data[616];
assign xnor2[617] = 1'b0 ^~ inbuffer_data[617];
assign xnor2[618] = 1'b0 ^~ inbuffer_data[618];
assign xnor2[619] = 1'b1 ^~ inbuffer_data[619];
assign xnor2[620] = 1'b1 ^~ inbuffer_data[620];
assign xnor2[621] = 1'b0 ^~ inbuffer_data[621];
assign xnor2[622] = 1'b1 ^~ inbuffer_data[622];
assign xnor2[623] = 1'b0 ^~ inbuffer_data[623];
assign xnor2[624] = 1'b1 ^~ inbuffer_data[624];
assign xnor2[625] = 1'b1 ^~ inbuffer_data[625];
assign xnor2[626] = 1'b0 ^~ inbuffer_data[626];
assign xnor2[627] = 1'b1 ^~ inbuffer_data[627];
assign xnor2[628] = 1'b1 ^~ inbuffer_data[628];
assign xnor2[629] = 1'b0 ^~ inbuffer_data[629];
assign xnor2[630] = 1'b1 ^~ inbuffer_data[630];
assign xnor2[631] = 1'b0 ^~ inbuffer_data[631];
assign xnor2[632] = 1'b0 ^~ inbuffer_data[632];
assign xnor2[633] = 1'b1 ^~ inbuffer_data[633];
assign xnor2[634] = 1'b1 ^~ inbuffer_data[634];
assign xnor2[635] = 1'b1 ^~ inbuffer_data[635];
assign xnor2[636] = 1'b1 ^~ inbuffer_data[636];
assign xnor2[637] = 1'b1 ^~ inbuffer_data[637];
assign xnor2[638] = 1'b1 ^~ inbuffer_data[638];
assign xnor2[639] = 1'b0 ^~ inbuffer_data[639];
assign xnor2[640] = 1'b1 ^~ inbuffer_data[640];
assign xnor2[641] = 1'b1 ^~ inbuffer_data[641];
assign xnor2[642] = 1'b0 ^~ inbuffer_data[642];
assign xnor2[643] = 1'b0 ^~ inbuffer_data[643];
assign xnor2[644] = 1'b0 ^~ inbuffer_data[644];
assign xnor2[645] = 1'b0 ^~ inbuffer_data[645];
assign xnor2[646] = 1'b0 ^~ inbuffer_data[646];
assign xnor2[647] = 1'b1 ^~ inbuffer_data[647];
assign xnor2[648] = 1'b0 ^~ inbuffer_data[648];
assign xnor2[649] = 1'b0 ^~ inbuffer_data[649];
assign xnor2[650] = 1'b0 ^~ inbuffer_data[650];
assign xnor2[651] = 1'b0 ^~ inbuffer_data[651];
assign xnor2[652] = 1'b1 ^~ inbuffer_data[652];
assign xnor2[653] = 1'b1 ^~ inbuffer_data[653];
assign xnor2[654] = 1'b1 ^~ inbuffer_data[654];
assign xnor2[655] = 1'b0 ^~ inbuffer_data[655];
assign xnor2[656] = 1'b0 ^~ inbuffer_data[656];
assign xnor2[657] = 1'b0 ^~ inbuffer_data[657];
assign xnor2[658] = 1'b0 ^~ inbuffer_data[658];
assign xnor2[659] = 1'b0 ^~ inbuffer_data[659];
assign xnor2[660] = 1'b0 ^~ inbuffer_data[660];
assign xnor2[661] = 1'b0 ^~ inbuffer_data[661];
assign xnor2[662] = 1'b1 ^~ inbuffer_data[662];
assign xnor2[663] = 1'b1 ^~ inbuffer_data[663];
assign xnor2[664] = 1'b1 ^~ inbuffer_data[664];
assign xnor2[665] = 1'b1 ^~ inbuffer_data[665];
assign xnor2[666] = 1'b1 ^~ inbuffer_data[666];
assign xnor2[667] = 1'b0 ^~ inbuffer_data[667];
assign xnor2[668] = 1'b0 ^~ inbuffer_data[668];
assign xnor2[669] = 1'b0 ^~ inbuffer_data[669];
assign xnor2[670] = 1'b1 ^~ inbuffer_data[670];
assign xnor2[671] = 1'b0 ^~ inbuffer_data[671];
assign xnor2[672] = 1'b0 ^~ inbuffer_data[672];
assign xnor2[673] = 1'b0 ^~ inbuffer_data[673];
assign xnor2[674] = 1'b0 ^~ inbuffer_data[674];
assign xnor2[675] = 1'b0 ^~ inbuffer_data[675];
assign xnor2[676] = 1'b0 ^~ inbuffer_data[676];
assign xnor2[677] = 1'b0 ^~ inbuffer_data[677];
assign xnor2[678] = 1'b0 ^~ inbuffer_data[678];
assign xnor2[679] = 1'b0 ^~ inbuffer_data[679];
assign xnor2[680] = 1'b0 ^~ inbuffer_data[680];
assign xnor2[681] = 1'b1 ^~ inbuffer_data[681];
assign xnor2[682] = 1'b0 ^~ inbuffer_data[682];
assign xnor2[683] = 1'b0 ^~ inbuffer_data[683];
assign xnor2[684] = 1'b0 ^~ inbuffer_data[684];
assign xnor2[685] = 1'b1 ^~ inbuffer_data[685];
assign xnor2[686] = 1'b1 ^~ inbuffer_data[686];
assign xnor2[687] = 1'b0 ^~ inbuffer_data[687];
assign xnor2[688] = 1'b1 ^~ inbuffer_data[688];
assign xnor2[689] = 1'b1 ^~ inbuffer_data[689];
assign xnor2[690] = 1'b1 ^~ inbuffer_data[690];
assign xnor2[691] = 1'b0 ^~ inbuffer_data[691];
assign xnor2[692] = 1'b0 ^~ inbuffer_data[692];
assign xnor2[693] = 1'b1 ^~ inbuffer_data[693];
assign xnor2[694] = 1'b0 ^~ inbuffer_data[694];
assign xnor2[695] = 1'b0 ^~ inbuffer_data[695];
assign xnor2[696] = 1'b0 ^~ inbuffer_data[696];
assign xnor2[697] = 1'b1 ^~ inbuffer_data[697];
assign xnor2[698] = 1'b1 ^~ inbuffer_data[698];
assign xnor2[699] = 1'b0 ^~ inbuffer_data[699];
assign xnor2[700] = 1'b1 ^~ inbuffer_data[700];
assign xnor2[701] = 1'b0 ^~ inbuffer_data[701];
assign xnor2[702] = 1'b0 ^~ inbuffer_data[702];
assign xnor2[703] = 1'b1 ^~ inbuffer_data[703];
assign xnor2[704] = 1'b1 ^~ inbuffer_data[704];
assign xnor2[705] = 1'b1 ^~ inbuffer_data[705];
assign xnor2[706] = 1'b0 ^~ inbuffer_data[706];
assign xnor2[707] = 1'b0 ^~ inbuffer_data[707];
assign xnor2[708] = 1'b0 ^~ inbuffer_data[708];
assign xnor2[709] = 1'b0 ^~ inbuffer_data[709];
assign xnor2[710] = 1'b0 ^~ inbuffer_data[710];
assign xnor2[711] = 1'b0 ^~ inbuffer_data[711];
assign xnor2[712] = 1'b0 ^~ inbuffer_data[712];
assign xnor2[713] = 1'b0 ^~ inbuffer_data[713];
assign xnor2[714] = 1'b0 ^~ inbuffer_data[714];
assign xnor2[715] = 1'b0 ^~ inbuffer_data[715];
assign xnor2[716] = 1'b0 ^~ inbuffer_data[716];
assign xnor2[717] = 1'b1 ^~ inbuffer_data[717];
assign xnor2[718] = 1'b0 ^~ inbuffer_data[718];
assign xnor2[719] = 1'b0 ^~ inbuffer_data[719];
assign xnor2[720] = 1'b0 ^~ inbuffer_data[720];
assign xnor2[721] = 1'b0 ^~ inbuffer_data[721];
assign xnor2[722] = 1'b0 ^~ inbuffer_data[722];
assign xnor2[723] = 1'b0 ^~ inbuffer_data[723];
assign xnor2[724] = 1'b0 ^~ inbuffer_data[724];
assign xnor2[725] = 1'b1 ^~ inbuffer_data[725];
assign xnor2[726] = 1'b1 ^~ inbuffer_data[726];
assign xnor2[727] = 1'b1 ^~ inbuffer_data[727];
assign xnor2[728] = 1'b0 ^~ inbuffer_data[728];
assign xnor2[729] = 1'b1 ^~ inbuffer_data[729];
assign xnor2[730] = 1'b0 ^~ inbuffer_data[730];
assign xnor2[731] = 1'b0 ^~ inbuffer_data[731];
assign xnor2[732] = 1'b0 ^~ inbuffer_data[732];
assign xnor2[733] = 1'b0 ^~ inbuffer_data[733];
assign xnor2[734] = 1'b1 ^~ inbuffer_data[734];
assign xnor2[735] = 1'b0 ^~ inbuffer_data[735];
assign xnor2[736] = 1'b1 ^~ inbuffer_data[736];
assign xnor2[737] = 1'b0 ^~ inbuffer_data[737];
assign xnor2[738] = 1'b0 ^~ inbuffer_data[738];
assign xnor2[739] = 1'b0 ^~ inbuffer_data[739];
assign xnor2[740] = 1'b1 ^~ inbuffer_data[740];
assign xnor2[741] = 1'b0 ^~ inbuffer_data[741];
assign xnor2[742] = 1'b0 ^~ inbuffer_data[742];
assign xnor2[743] = 1'b0 ^~ inbuffer_data[743];
assign xnor2[744] = 1'b0 ^~ inbuffer_data[744];
assign xnor2[745] = 1'b0 ^~ inbuffer_data[745];
assign xnor2[746] = 1'b0 ^~ inbuffer_data[746];
assign xnor2[747] = 1'b0 ^~ inbuffer_data[747];
assign xnor2[748] = 1'b0 ^~ inbuffer_data[748];
assign xnor2[749] = 1'b0 ^~ inbuffer_data[749];
assign xnor2[750] = 1'b1 ^~ inbuffer_data[750];
assign xnor2[751] = 1'b0 ^~ inbuffer_data[751];
assign xnor2[752] = 1'b1 ^~ inbuffer_data[752];
assign xnor2[753] = 1'b0 ^~ inbuffer_data[753];
assign xnor2[754] = 1'b0 ^~ inbuffer_data[754];
assign xnor2[755] = 1'b0 ^~ inbuffer_data[755];
assign xnor2[756] = 1'b0 ^~ inbuffer_data[756];
assign xnor2[757] = 1'b0 ^~ inbuffer_data[757];
assign xnor2[758] = 1'b1 ^~ inbuffer_data[758];
assign xnor2[759] = 1'b1 ^~ inbuffer_data[759];
assign xnor2[760] = 1'b0 ^~ inbuffer_data[760];
assign xnor2[761] = 1'b0 ^~ inbuffer_data[761];
assign xnor2[762] = 1'b0 ^~ inbuffer_data[762];
assign xnor2[763] = 1'b0 ^~ inbuffer_data[763];
assign xnor2[764] = 1'b0 ^~ inbuffer_data[764];
assign xnor2[765] = 1'b0 ^~ inbuffer_data[765];
assign xnor2[766] = 1'b0 ^~ inbuffer_data[766];
assign xnor2[767] = 1'b0 ^~ inbuffer_data[767];
assign xnor2[768] = 1'b0 ^~ inbuffer_data[768];
assign xnor2[769] = 1'b0 ^~ inbuffer_data[769];
assign xnor2[770] = 1'b1 ^~ inbuffer_data[770];
assign xnor2[771] = 1'b0 ^~ inbuffer_data[771];
assign xnor2[772] = 1'b1 ^~ inbuffer_data[772];
assign xnor2[773] = 1'b1 ^~ inbuffer_data[773];
assign xnor2[774] = 1'b0 ^~ inbuffer_data[774];
assign xnor2[775] = 1'b0 ^~ inbuffer_data[775];
assign xnor2[776] = 1'b1 ^~ inbuffer_data[776];
assign xnor2[777] = 1'b1 ^~ inbuffer_data[777];
assign xnor2[778] = 1'b0 ^~ inbuffer_data[778];
assign xnor2[779] = 1'b0 ^~ inbuffer_data[779];
assign xnor2[780] = 1'b0 ^~ inbuffer_data[780];
assign xnor2[781] = 1'b0 ^~ inbuffer_data[781];
assign xnor2[782] = 1'b0 ^~ inbuffer_data[782];
assign xnor2[783] = 1'b1 ^~ inbuffer_data[783];
assign xnor3[0] = 1'b0 ^~ inbuffer_data[0];
assign xnor3[1] = 1'b0 ^~ inbuffer_data[1];
assign xnor3[2] = 1'b1 ^~ inbuffer_data[2];
assign xnor3[3] = 1'b1 ^~ inbuffer_data[3];
assign xnor3[4] = 1'b0 ^~ inbuffer_data[4];
assign xnor3[5] = 1'b1 ^~ inbuffer_data[5];
assign xnor3[6] = 1'b1 ^~ inbuffer_data[6];
assign xnor3[7] = 1'b0 ^~ inbuffer_data[7];
assign xnor3[8] = 1'b0 ^~ inbuffer_data[8];
assign xnor3[9] = 1'b0 ^~ inbuffer_data[9];
assign xnor3[10] = 1'b0 ^~ inbuffer_data[10];
assign xnor3[11] = 1'b0 ^~ inbuffer_data[11];
assign xnor3[12] = 1'b1 ^~ inbuffer_data[12];
assign xnor3[13] = 1'b0 ^~ inbuffer_data[13];
assign xnor3[14] = 1'b0 ^~ inbuffer_data[14];
assign xnor3[15] = 1'b0 ^~ inbuffer_data[15];
assign xnor3[16] = 1'b1 ^~ inbuffer_data[16];
assign xnor3[17] = 1'b0 ^~ inbuffer_data[17];
assign xnor3[18] = 1'b1 ^~ inbuffer_data[18];
assign xnor3[19] = 1'b0 ^~ inbuffer_data[19];
assign xnor3[20] = 1'b0 ^~ inbuffer_data[20];
assign xnor3[21] = 1'b1 ^~ inbuffer_data[21];
assign xnor3[22] = 1'b0 ^~ inbuffer_data[22];
assign xnor3[23] = 1'b1 ^~ inbuffer_data[23];
assign xnor3[24] = 1'b1 ^~ inbuffer_data[24];
assign xnor3[25] = 1'b0 ^~ inbuffer_data[25];
assign xnor3[26] = 1'b0 ^~ inbuffer_data[26];
assign xnor3[27] = 1'b1 ^~ inbuffer_data[27];
assign xnor3[28] = 1'b0 ^~ inbuffer_data[28];
assign xnor3[29] = 1'b0 ^~ inbuffer_data[29];
assign xnor3[30] = 1'b0 ^~ inbuffer_data[30];
assign xnor3[31] = 1'b0 ^~ inbuffer_data[31];
assign xnor3[32] = 1'b0 ^~ inbuffer_data[32];
assign xnor3[33] = 1'b0 ^~ inbuffer_data[33];
assign xnor3[34] = 1'b1 ^~ inbuffer_data[34];
assign xnor3[35] = 1'b1 ^~ inbuffer_data[35];
assign xnor3[36] = 1'b0 ^~ inbuffer_data[36];
assign xnor3[37] = 1'b0 ^~ inbuffer_data[37];
assign xnor3[38] = 1'b1 ^~ inbuffer_data[38];
assign xnor3[39] = 1'b1 ^~ inbuffer_data[39];
assign xnor3[40] = 1'b0 ^~ inbuffer_data[40];
assign xnor3[41] = 1'b1 ^~ inbuffer_data[41];
assign xnor3[42] = 1'b0 ^~ inbuffer_data[42];
assign xnor3[43] = 1'b1 ^~ inbuffer_data[43];
assign xnor3[44] = 1'b0 ^~ inbuffer_data[44];
assign xnor3[45] = 1'b0 ^~ inbuffer_data[45];
assign xnor3[46] = 1'b1 ^~ inbuffer_data[46];
assign xnor3[47] = 1'b1 ^~ inbuffer_data[47];
assign xnor3[48] = 1'b0 ^~ inbuffer_data[48];
assign xnor3[49] = 1'b1 ^~ inbuffer_data[49];
assign xnor3[50] = 1'b1 ^~ inbuffer_data[50];
assign xnor3[51] = 1'b0 ^~ inbuffer_data[51];
assign xnor3[52] = 1'b0 ^~ inbuffer_data[52];
assign xnor3[53] = 1'b0 ^~ inbuffer_data[53];
assign xnor3[54] = 1'b0 ^~ inbuffer_data[54];
assign xnor3[55] = 1'b0 ^~ inbuffer_data[55];
assign xnor3[56] = 1'b0 ^~ inbuffer_data[56];
assign xnor3[57] = 1'b0 ^~ inbuffer_data[57];
assign xnor3[58] = 1'b1 ^~ inbuffer_data[58];
assign xnor3[59] = 1'b1 ^~ inbuffer_data[59];
assign xnor3[60] = 1'b0 ^~ inbuffer_data[60];
assign xnor3[61] = 1'b0 ^~ inbuffer_data[61];
assign xnor3[62] = 1'b0 ^~ inbuffer_data[62];
assign xnor3[63] = 1'b0 ^~ inbuffer_data[63];
assign xnor3[64] = 1'b1 ^~ inbuffer_data[64];
assign xnor3[65] = 1'b0 ^~ inbuffer_data[65];
assign xnor3[66] = 1'b0 ^~ inbuffer_data[66];
assign xnor3[67] = 1'b1 ^~ inbuffer_data[67];
assign xnor3[68] = 1'b0 ^~ inbuffer_data[68];
assign xnor3[69] = 1'b0 ^~ inbuffer_data[69];
assign xnor3[70] = 1'b0 ^~ inbuffer_data[70];
assign xnor3[71] = 1'b1 ^~ inbuffer_data[71];
assign xnor3[72] = 1'b1 ^~ inbuffer_data[72];
assign xnor3[73] = 1'b0 ^~ inbuffer_data[73];
assign xnor3[74] = 1'b0 ^~ inbuffer_data[74];
assign xnor3[75] = 1'b1 ^~ inbuffer_data[75];
assign xnor3[76] = 1'b1 ^~ inbuffer_data[76];
assign xnor3[77] = 1'b0 ^~ inbuffer_data[77];
assign xnor3[78] = 1'b0 ^~ inbuffer_data[78];
assign xnor3[79] = 1'b1 ^~ inbuffer_data[79];
assign xnor3[80] = 1'b0 ^~ inbuffer_data[80];
assign xnor3[81] = 1'b0 ^~ inbuffer_data[81];
assign xnor3[82] = 1'b1 ^~ inbuffer_data[82];
assign xnor3[83] = 1'b0 ^~ inbuffer_data[83];
assign xnor3[84] = 1'b0 ^~ inbuffer_data[84];
assign xnor3[85] = 1'b0 ^~ inbuffer_data[85];
assign xnor3[86] = 1'b0 ^~ inbuffer_data[86];
assign xnor3[87] = 1'b1 ^~ inbuffer_data[87];
assign xnor3[88] = 1'b0 ^~ inbuffer_data[88];
assign xnor3[89] = 1'b1 ^~ inbuffer_data[89];
assign xnor3[90] = 1'b0 ^~ inbuffer_data[90];
assign xnor3[91] = 1'b0 ^~ inbuffer_data[91];
assign xnor3[92] = 1'b0 ^~ inbuffer_data[92];
assign xnor3[93] = 1'b1 ^~ inbuffer_data[93];
assign xnor3[94] = 1'b0 ^~ inbuffer_data[94];
assign xnor3[95] = 1'b1 ^~ inbuffer_data[95];
assign xnor3[96] = 1'b1 ^~ inbuffer_data[96];
assign xnor3[97] = 1'b1 ^~ inbuffer_data[97];
assign xnor3[98] = 1'b1 ^~ inbuffer_data[98];
assign xnor3[99] = 1'b1 ^~ inbuffer_data[99];
assign xnor3[100] = 1'b1 ^~ inbuffer_data[100];
assign xnor3[101] = 1'b1 ^~ inbuffer_data[101];
assign xnor3[102] = 1'b1 ^~ inbuffer_data[102];
assign xnor3[103] = 1'b1 ^~ inbuffer_data[103];
assign xnor3[104] = 1'b0 ^~ inbuffer_data[104];
assign xnor3[105] = 1'b0 ^~ inbuffer_data[105];
assign xnor3[106] = 1'b0 ^~ inbuffer_data[106];
assign xnor3[107] = 1'b0 ^~ inbuffer_data[107];
assign xnor3[108] = 1'b0 ^~ inbuffer_data[108];
assign xnor3[109] = 1'b0 ^~ inbuffer_data[109];
assign xnor3[110] = 1'b0 ^~ inbuffer_data[110];
assign xnor3[111] = 1'b0 ^~ inbuffer_data[111];
assign xnor3[112] = 1'b0 ^~ inbuffer_data[112];
assign xnor3[113] = 1'b1 ^~ inbuffer_data[113];
assign xnor3[114] = 1'b0 ^~ inbuffer_data[114];
assign xnor3[115] = 1'b0 ^~ inbuffer_data[115];
assign xnor3[116] = 1'b1 ^~ inbuffer_data[116];
assign xnor3[117] = 1'b1 ^~ inbuffer_data[117];
assign xnor3[118] = 1'b1 ^~ inbuffer_data[118];
assign xnor3[119] = 1'b1 ^~ inbuffer_data[119];
assign xnor3[120] = 1'b1 ^~ inbuffer_data[120];
assign xnor3[121] = 1'b1 ^~ inbuffer_data[121];
assign xnor3[122] = 1'b1 ^~ inbuffer_data[122];
assign xnor3[123] = 1'b1 ^~ inbuffer_data[123];
assign xnor3[124] = 1'b1 ^~ inbuffer_data[124];
assign xnor3[125] = 1'b1 ^~ inbuffer_data[125];
assign xnor3[126] = 1'b1 ^~ inbuffer_data[126];
assign xnor3[127] = 1'b1 ^~ inbuffer_data[127];
assign xnor3[128] = 1'b1 ^~ inbuffer_data[128];
assign xnor3[129] = 1'b1 ^~ inbuffer_data[129];
assign xnor3[130] = 1'b1 ^~ inbuffer_data[130];
assign xnor3[131] = 1'b1 ^~ inbuffer_data[131];
assign xnor3[132] = 1'b1 ^~ inbuffer_data[132];
assign xnor3[133] = 1'b0 ^~ inbuffer_data[133];
assign xnor3[134] = 1'b0 ^~ inbuffer_data[134];
assign xnor3[135] = 1'b0 ^~ inbuffer_data[135];
assign xnor3[136] = 1'b1 ^~ inbuffer_data[136];
assign xnor3[137] = 1'b1 ^~ inbuffer_data[137];
assign xnor3[138] = 1'b1 ^~ inbuffer_data[138];
assign xnor3[139] = 1'b1 ^~ inbuffer_data[139];
assign xnor3[140] = 1'b0 ^~ inbuffer_data[140];
assign xnor3[141] = 1'b0 ^~ inbuffer_data[141];
assign xnor3[142] = 1'b0 ^~ inbuffer_data[142];
assign xnor3[143] = 1'b1 ^~ inbuffer_data[143];
assign xnor3[144] = 1'b1 ^~ inbuffer_data[144];
assign xnor3[145] = 1'b1 ^~ inbuffer_data[145];
assign xnor3[146] = 1'b1 ^~ inbuffer_data[146];
assign xnor3[147] = 1'b1 ^~ inbuffer_data[147];
assign xnor3[148] = 1'b1 ^~ inbuffer_data[148];
assign xnor3[149] = 1'b1 ^~ inbuffer_data[149];
assign xnor3[150] = 1'b1 ^~ inbuffer_data[150];
assign xnor3[151] = 1'b1 ^~ inbuffer_data[151];
assign xnor3[152] = 1'b1 ^~ inbuffer_data[152];
assign xnor3[153] = 1'b0 ^~ inbuffer_data[153];
assign xnor3[154] = 1'b0 ^~ inbuffer_data[154];
assign xnor3[155] = 1'b1 ^~ inbuffer_data[155];
assign xnor3[156] = 1'b1 ^~ inbuffer_data[156];
assign xnor3[157] = 1'b1 ^~ inbuffer_data[157];
assign xnor3[158] = 1'b1 ^~ inbuffer_data[158];
assign xnor3[159] = 1'b1 ^~ inbuffer_data[159];
assign xnor3[160] = 1'b0 ^~ inbuffer_data[160];
assign xnor3[161] = 1'b0 ^~ inbuffer_data[161];
assign xnor3[162] = 1'b0 ^~ inbuffer_data[162];
assign xnor3[163] = 1'b0 ^~ inbuffer_data[163];
assign xnor3[164] = 1'b1 ^~ inbuffer_data[164];
assign xnor3[165] = 1'b1 ^~ inbuffer_data[165];
assign xnor3[166] = 1'b1 ^~ inbuffer_data[166];
assign xnor3[167] = 1'b0 ^~ inbuffer_data[167];
assign xnor3[168] = 1'b1 ^~ inbuffer_data[168];
assign xnor3[169] = 1'b0 ^~ inbuffer_data[169];
assign xnor3[170] = 1'b0 ^~ inbuffer_data[170];
assign xnor3[171] = 1'b1 ^~ inbuffer_data[171];
assign xnor3[172] = 1'b1 ^~ inbuffer_data[172];
assign xnor3[173] = 1'b1 ^~ inbuffer_data[173];
assign xnor3[174] = 1'b1 ^~ inbuffer_data[174];
assign xnor3[175] = 1'b1 ^~ inbuffer_data[175];
assign xnor3[176] = 1'b1 ^~ inbuffer_data[176];
assign xnor3[177] = 1'b1 ^~ inbuffer_data[177];
assign xnor3[178] = 1'b1 ^~ inbuffer_data[178];
assign xnor3[179] = 1'b0 ^~ inbuffer_data[179];
assign xnor3[180] = 1'b1 ^~ inbuffer_data[180];
assign xnor3[181] = 1'b1 ^~ inbuffer_data[181];
assign xnor3[182] = 1'b1 ^~ inbuffer_data[182];
assign xnor3[183] = 1'b1 ^~ inbuffer_data[183];
assign xnor3[184] = 1'b1 ^~ inbuffer_data[184];
assign xnor3[185] = 1'b0 ^~ inbuffer_data[185];
assign xnor3[186] = 1'b1 ^~ inbuffer_data[186];
assign xnor3[187] = 1'b0 ^~ inbuffer_data[187];
assign xnor3[188] = 1'b1 ^~ inbuffer_data[188];
assign xnor3[189] = 1'b1 ^~ inbuffer_data[189];
assign xnor3[190] = 1'b0 ^~ inbuffer_data[190];
assign xnor3[191] = 1'b0 ^~ inbuffer_data[191];
assign xnor3[192] = 1'b0 ^~ inbuffer_data[192];
assign xnor3[193] = 1'b0 ^~ inbuffer_data[193];
assign xnor3[194] = 1'b0 ^~ inbuffer_data[194];
assign xnor3[195] = 1'b0 ^~ inbuffer_data[195];
assign xnor3[196] = 1'b0 ^~ inbuffer_data[196];
assign xnor3[197] = 1'b0 ^~ inbuffer_data[197];
assign xnor3[198] = 1'b0 ^~ inbuffer_data[198];
assign xnor3[199] = 1'b1 ^~ inbuffer_data[199];
assign xnor3[200] = 1'b1 ^~ inbuffer_data[200];
assign xnor3[201] = 1'b1 ^~ inbuffer_data[201];
assign xnor3[202] = 1'b1 ^~ inbuffer_data[202];
assign xnor3[203] = 1'b1 ^~ inbuffer_data[203];
assign xnor3[204] = 1'b1 ^~ inbuffer_data[204];
assign xnor3[205] = 1'b1 ^~ inbuffer_data[205];
assign xnor3[206] = 1'b0 ^~ inbuffer_data[206];
assign xnor3[207] = 1'b1 ^~ inbuffer_data[207];
assign xnor3[208] = 1'b1 ^~ inbuffer_data[208];
assign xnor3[209] = 1'b0 ^~ inbuffer_data[209];
assign xnor3[210] = 1'b1 ^~ inbuffer_data[210];
assign xnor3[211] = 1'b1 ^~ inbuffer_data[211];
assign xnor3[212] = 1'b0 ^~ inbuffer_data[212];
assign xnor3[213] = 1'b0 ^~ inbuffer_data[213];
assign xnor3[214] = 1'b1 ^~ inbuffer_data[214];
assign xnor3[215] = 1'b1 ^~ inbuffer_data[215];
assign xnor3[216] = 1'b0 ^~ inbuffer_data[216];
assign xnor3[217] = 1'b1 ^~ inbuffer_data[217];
assign xnor3[218] = 1'b0 ^~ inbuffer_data[218];
assign xnor3[219] = 1'b0 ^~ inbuffer_data[219];
assign xnor3[220] = 1'b0 ^~ inbuffer_data[220];
assign xnor3[221] = 1'b0 ^~ inbuffer_data[221];
assign xnor3[222] = 1'b1 ^~ inbuffer_data[222];
assign xnor3[223] = 1'b0 ^~ inbuffer_data[223];
assign xnor3[224] = 1'b1 ^~ inbuffer_data[224];
assign xnor3[225] = 1'b0 ^~ inbuffer_data[225];
assign xnor3[226] = 1'b0 ^~ inbuffer_data[226];
assign xnor3[227] = 1'b0 ^~ inbuffer_data[227];
assign xnor3[228] = 1'b1 ^~ inbuffer_data[228];
assign xnor3[229] = 1'b1 ^~ inbuffer_data[229];
assign xnor3[230] = 1'b1 ^~ inbuffer_data[230];
assign xnor3[231] = 1'b1 ^~ inbuffer_data[231];
assign xnor3[232] = 1'b1 ^~ inbuffer_data[232];
assign xnor3[233] = 1'b1 ^~ inbuffer_data[233];
assign xnor3[234] = 1'b1 ^~ inbuffer_data[234];
assign xnor3[235] = 1'b0 ^~ inbuffer_data[235];
assign xnor3[236] = 1'b1 ^~ inbuffer_data[236];
assign xnor3[237] = 1'b1 ^~ inbuffer_data[237];
assign xnor3[238] = 1'b1 ^~ inbuffer_data[238];
assign xnor3[239] = 1'b1 ^~ inbuffer_data[239];
assign xnor3[240] = 1'b1 ^~ inbuffer_data[240];
assign xnor3[241] = 1'b1 ^~ inbuffer_data[241];
assign xnor3[242] = 1'b1 ^~ inbuffer_data[242];
assign xnor3[243] = 1'b1 ^~ inbuffer_data[243];
assign xnor3[244] = 1'b1 ^~ inbuffer_data[244];
assign xnor3[245] = 1'b1 ^~ inbuffer_data[245];
assign xnor3[246] = 1'b0 ^~ inbuffer_data[246];
assign xnor3[247] = 1'b0 ^~ inbuffer_data[247];
assign xnor3[248] = 1'b0 ^~ inbuffer_data[248];
assign xnor3[249] = 1'b0 ^~ inbuffer_data[249];
assign xnor3[250] = 1'b0 ^~ inbuffer_data[250];
assign xnor3[251] = 1'b0 ^~ inbuffer_data[251];
assign xnor3[252] = 1'b0 ^~ inbuffer_data[252];
assign xnor3[253] = 1'b0 ^~ inbuffer_data[253];
assign xnor3[254] = 1'b1 ^~ inbuffer_data[254];
assign xnor3[255] = 1'b1 ^~ inbuffer_data[255];
assign xnor3[256] = 1'b1 ^~ inbuffer_data[256];
assign xnor3[257] = 1'b1 ^~ inbuffer_data[257];
assign xnor3[258] = 1'b0 ^~ inbuffer_data[258];
assign xnor3[259] = 1'b1 ^~ inbuffer_data[259];
assign xnor3[260] = 1'b0 ^~ inbuffer_data[260];
assign xnor3[261] = 1'b0 ^~ inbuffer_data[261];
assign xnor3[262] = 1'b0 ^~ inbuffer_data[262];
assign xnor3[263] = 1'b0 ^~ inbuffer_data[263];
assign xnor3[264] = 1'b0 ^~ inbuffer_data[264];
assign xnor3[265] = 1'b0 ^~ inbuffer_data[265];
assign xnor3[266] = 1'b1 ^~ inbuffer_data[266];
assign xnor3[267] = 1'b1 ^~ inbuffer_data[267];
assign xnor3[268] = 1'b0 ^~ inbuffer_data[268];
assign xnor3[269] = 1'b0 ^~ inbuffer_data[269];
assign xnor3[270] = 1'b1 ^~ inbuffer_data[270];
assign xnor3[271] = 1'b1 ^~ inbuffer_data[271];
assign xnor3[272] = 1'b1 ^~ inbuffer_data[272];
assign xnor3[273] = 1'b1 ^~ inbuffer_data[273];
assign xnor3[274] = 1'b1 ^~ inbuffer_data[274];
assign xnor3[275] = 1'b0 ^~ inbuffer_data[275];
assign xnor3[276] = 1'b0 ^~ inbuffer_data[276];
assign xnor3[277] = 1'b0 ^~ inbuffer_data[277];
assign xnor3[278] = 1'b0 ^~ inbuffer_data[278];
assign xnor3[279] = 1'b1 ^~ inbuffer_data[279];
assign xnor3[280] = 1'b0 ^~ inbuffer_data[280];
assign xnor3[281] = 1'b0 ^~ inbuffer_data[281];
assign xnor3[282] = 1'b1 ^~ inbuffer_data[282];
assign xnor3[283] = 1'b1 ^~ inbuffer_data[283];
assign xnor3[284] = 1'b1 ^~ inbuffer_data[284];
assign xnor3[285] = 1'b1 ^~ inbuffer_data[285];
assign xnor3[286] = 1'b0 ^~ inbuffer_data[286];
assign xnor3[287] = 1'b0 ^~ inbuffer_data[287];
assign xnor3[288] = 1'b0 ^~ inbuffer_data[288];
assign xnor3[289] = 1'b0 ^~ inbuffer_data[289];
assign xnor3[290] = 1'b0 ^~ inbuffer_data[290];
assign xnor3[291] = 1'b0 ^~ inbuffer_data[291];
assign xnor3[292] = 1'b0 ^~ inbuffer_data[292];
assign xnor3[293] = 1'b0 ^~ inbuffer_data[293];
assign xnor3[294] = 1'b1 ^~ inbuffer_data[294];
assign xnor3[295] = 1'b1 ^~ inbuffer_data[295];
assign xnor3[296] = 1'b1 ^~ inbuffer_data[296];
assign xnor3[297] = 1'b1 ^~ inbuffer_data[297];
assign xnor3[298] = 1'b1 ^~ inbuffer_data[298];
assign xnor3[299] = 1'b1 ^~ inbuffer_data[299];
assign xnor3[300] = 1'b1 ^~ inbuffer_data[300];
assign xnor3[301] = 1'b1 ^~ inbuffer_data[301];
assign xnor3[302] = 1'b1 ^~ inbuffer_data[302];
assign xnor3[303] = 1'b0 ^~ inbuffer_data[303];
assign xnor3[304] = 1'b0 ^~ inbuffer_data[304];
assign xnor3[305] = 1'b0 ^~ inbuffer_data[305];
assign xnor3[306] = 1'b0 ^~ inbuffer_data[306];
assign xnor3[307] = 1'b0 ^~ inbuffer_data[307];
assign xnor3[308] = 1'b0 ^~ inbuffer_data[308];
assign xnor3[309] = 1'b0 ^~ inbuffer_data[309];
assign xnor3[310] = 1'b1 ^~ inbuffer_data[310];
assign xnor3[311] = 1'b1 ^~ inbuffer_data[311];
assign xnor3[312] = 1'b1 ^~ inbuffer_data[312];
assign xnor3[313] = 1'b0 ^~ inbuffer_data[313];
assign xnor3[314] = 1'b0 ^~ inbuffer_data[314];
assign xnor3[315] = 1'b0 ^~ inbuffer_data[315];
assign xnor3[316] = 1'b0 ^~ inbuffer_data[316];
assign xnor3[317] = 1'b0 ^~ inbuffer_data[317];
assign xnor3[318] = 1'b0 ^~ inbuffer_data[318];
assign xnor3[319] = 1'b0 ^~ inbuffer_data[319];
assign xnor3[320] = 1'b0 ^~ inbuffer_data[320];
assign xnor3[321] = 1'b1 ^~ inbuffer_data[321];
assign xnor3[322] = 1'b1 ^~ inbuffer_data[322];
assign xnor3[323] = 1'b1 ^~ inbuffer_data[323];
assign xnor3[324] = 1'b0 ^~ inbuffer_data[324];
assign xnor3[325] = 1'b1 ^~ inbuffer_data[325];
assign xnor3[326] = 1'b1 ^~ inbuffer_data[326];
assign xnor3[327] = 1'b1 ^~ inbuffer_data[327];
assign xnor3[328] = 1'b1 ^~ inbuffer_data[328];
assign xnor3[329] = 1'b0 ^~ inbuffer_data[329];
assign xnor3[330] = 1'b1 ^~ inbuffer_data[330];
assign xnor3[331] = 1'b0 ^~ inbuffer_data[331];
assign xnor3[332] = 1'b0 ^~ inbuffer_data[332];
assign xnor3[333] = 1'b0 ^~ inbuffer_data[333];
assign xnor3[334] = 1'b1 ^~ inbuffer_data[334];
assign xnor3[335] = 1'b0 ^~ inbuffer_data[335];
assign xnor3[336] = 1'b1 ^~ inbuffer_data[336];
assign xnor3[337] = 1'b0 ^~ inbuffer_data[337];
assign xnor3[338] = 1'b0 ^~ inbuffer_data[338];
assign xnor3[339] = 1'b0 ^~ inbuffer_data[339];
assign xnor3[340] = 1'b0 ^~ inbuffer_data[340];
assign xnor3[341] = 1'b0 ^~ inbuffer_data[341];
assign xnor3[342] = 1'b0 ^~ inbuffer_data[342];
assign xnor3[343] = 1'b0 ^~ inbuffer_data[343];
assign xnor3[344] = 1'b0 ^~ inbuffer_data[344];
assign xnor3[345] = 1'b0 ^~ inbuffer_data[345];
assign xnor3[346] = 1'b1 ^~ inbuffer_data[346];
assign xnor3[347] = 1'b0 ^~ inbuffer_data[347];
assign xnor3[348] = 1'b1 ^~ inbuffer_data[348];
assign xnor3[349] = 1'b1 ^~ inbuffer_data[349];
assign xnor3[350] = 1'b1 ^~ inbuffer_data[350];
assign xnor3[351] = 1'b1 ^~ inbuffer_data[351];
assign xnor3[352] = 1'b1 ^~ inbuffer_data[352];
assign xnor3[353] = 1'b1 ^~ inbuffer_data[353];
assign xnor3[354] = 1'b1 ^~ inbuffer_data[354];
assign xnor3[355] = 1'b1 ^~ inbuffer_data[355];
assign xnor3[356] = 1'b0 ^~ inbuffer_data[356];
assign xnor3[357] = 1'b0 ^~ inbuffer_data[357];
assign xnor3[358] = 1'b0 ^~ inbuffer_data[358];
assign xnor3[359] = 1'b0 ^~ inbuffer_data[359];
assign xnor3[360] = 1'b0 ^~ inbuffer_data[360];
assign xnor3[361] = 1'b0 ^~ inbuffer_data[361];
assign xnor3[362] = 1'b0 ^~ inbuffer_data[362];
assign xnor3[363] = 1'b0 ^~ inbuffer_data[363];
assign xnor3[364] = 1'b0 ^~ inbuffer_data[364];
assign xnor3[365] = 1'b1 ^~ inbuffer_data[365];
assign xnor3[366] = 1'b1 ^~ inbuffer_data[366];
assign xnor3[367] = 1'b0 ^~ inbuffer_data[367];
assign xnor3[368] = 1'b0 ^~ inbuffer_data[368];
assign xnor3[369] = 1'b0 ^~ inbuffer_data[369];
assign xnor3[370] = 1'b0 ^~ inbuffer_data[370];
assign xnor3[371] = 1'b0 ^~ inbuffer_data[371];
assign xnor3[372] = 1'b0 ^~ inbuffer_data[372];
assign xnor3[373] = 1'b0 ^~ inbuffer_data[373];
assign xnor3[374] = 1'b0 ^~ inbuffer_data[374];
assign xnor3[375] = 1'b1 ^~ inbuffer_data[375];
assign xnor3[376] = 1'b0 ^~ inbuffer_data[376];
assign xnor3[377] = 1'b1 ^~ inbuffer_data[377];
assign xnor3[378] = 1'b1 ^~ inbuffer_data[378];
assign xnor3[379] = 1'b1 ^~ inbuffer_data[379];
assign xnor3[380] = 1'b1 ^~ inbuffer_data[380];
assign xnor3[381] = 1'b1 ^~ inbuffer_data[381];
assign xnor3[382] = 1'b0 ^~ inbuffer_data[382];
assign xnor3[383] = 1'b0 ^~ inbuffer_data[383];
assign xnor3[384] = 1'b0 ^~ inbuffer_data[384];
assign xnor3[385] = 1'b0 ^~ inbuffer_data[385];
assign xnor3[386] = 1'b0 ^~ inbuffer_data[386];
assign xnor3[387] = 1'b0 ^~ inbuffer_data[387];
assign xnor3[388] = 1'b1 ^~ inbuffer_data[388];
assign xnor3[389] = 1'b0 ^~ inbuffer_data[389];
assign xnor3[390] = 1'b0 ^~ inbuffer_data[390];
assign xnor3[391] = 1'b1 ^~ inbuffer_data[391];
assign xnor3[392] = 1'b1 ^~ inbuffer_data[392];
assign xnor3[393] = 1'b0 ^~ inbuffer_data[393];
assign xnor3[394] = 1'b0 ^~ inbuffer_data[394];
assign xnor3[395] = 1'b1 ^~ inbuffer_data[395];
assign xnor3[396] = 1'b0 ^~ inbuffer_data[396];
assign xnor3[397] = 1'b0 ^~ inbuffer_data[397];
assign xnor3[398] = 1'b0 ^~ inbuffer_data[398];
assign xnor3[399] = 1'b0 ^~ inbuffer_data[399];
assign xnor3[400] = 1'b0 ^~ inbuffer_data[400];
assign xnor3[401] = 1'b1 ^~ inbuffer_data[401];
assign xnor3[402] = 1'b0 ^~ inbuffer_data[402];
assign xnor3[403] = 1'b1 ^~ inbuffer_data[403];
assign xnor3[404] = 1'b1 ^~ inbuffer_data[404];
assign xnor3[405] = 1'b0 ^~ inbuffer_data[405];
assign xnor3[406] = 1'b1 ^~ inbuffer_data[406];
assign xnor3[407] = 1'b1 ^~ inbuffer_data[407];
assign xnor3[408] = 1'b0 ^~ inbuffer_data[408];
assign xnor3[409] = 1'b1 ^~ inbuffer_data[409];
assign xnor3[410] = 1'b0 ^~ inbuffer_data[410];
assign xnor3[411] = 1'b0 ^~ inbuffer_data[411];
assign xnor3[412] = 1'b0 ^~ inbuffer_data[412];
assign xnor3[413] = 1'b1 ^~ inbuffer_data[413];
assign xnor3[414] = 1'b0 ^~ inbuffer_data[414];
assign xnor3[415] = 1'b0 ^~ inbuffer_data[415];
assign xnor3[416] = 1'b0 ^~ inbuffer_data[416];
assign xnor3[417] = 1'b1 ^~ inbuffer_data[417];
assign xnor3[418] = 1'b1 ^~ inbuffer_data[418];
assign xnor3[419] = 1'b1 ^~ inbuffer_data[419];
assign xnor3[420] = 1'b0 ^~ inbuffer_data[420];
assign xnor3[421] = 1'b0 ^~ inbuffer_data[421];
assign xnor3[422] = 1'b0 ^~ inbuffer_data[422];
assign xnor3[423] = 1'b1 ^~ inbuffer_data[423];
assign xnor3[424] = 1'b1 ^~ inbuffer_data[424];
assign xnor3[425] = 1'b1 ^~ inbuffer_data[425];
assign xnor3[426] = 1'b0 ^~ inbuffer_data[426];
assign xnor3[427] = 1'b0 ^~ inbuffer_data[427];
assign xnor3[428] = 1'b0 ^~ inbuffer_data[428];
assign xnor3[429] = 1'b0 ^~ inbuffer_data[429];
assign xnor3[430] = 1'b0 ^~ inbuffer_data[430];
assign xnor3[431] = 1'b1 ^~ inbuffer_data[431];
assign xnor3[432] = 1'b1 ^~ inbuffer_data[432];
assign xnor3[433] = 1'b0 ^~ inbuffer_data[433];
assign xnor3[434] = 1'b1 ^~ inbuffer_data[434];
assign xnor3[435] = 1'b1 ^~ inbuffer_data[435];
assign xnor3[436] = 1'b0 ^~ inbuffer_data[436];
assign xnor3[437] = 1'b1 ^~ inbuffer_data[437];
assign xnor3[438] = 1'b0 ^~ inbuffer_data[438];
assign xnor3[439] = 1'b1 ^~ inbuffer_data[439];
assign xnor3[440] = 1'b1 ^~ inbuffer_data[440];
assign xnor3[441] = 1'b0 ^~ inbuffer_data[441];
assign xnor3[442] = 1'b1 ^~ inbuffer_data[442];
assign xnor3[443] = 1'b1 ^~ inbuffer_data[443];
assign xnor3[444] = 1'b0 ^~ inbuffer_data[444];
assign xnor3[445] = 1'b0 ^~ inbuffer_data[445];
assign xnor3[446] = 1'b1 ^~ inbuffer_data[446];
assign xnor3[447] = 1'b0 ^~ inbuffer_data[447];
assign xnor3[448] = 1'b0 ^~ inbuffer_data[448];
assign xnor3[449] = 1'b0 ^~ inbuffer_data[449];
assign xnor3[450] = 1'b1 ^~ inbuffer_data[450];
assign xnor3[451] = 1'b0 ^~ inbuffer_data[451];
assign xnor3[452] = 1'b1 ^~ inbuffer_data[452];
assign xnor3[453] = 1'b1 ^~ inbuffer_data[453];
assign xnor3[454] = 1'b0 ^~ inbuffer_data[454];
assign xnor3[455] = 1'b0 ^~ inbuffer_data[455];
assign xnor3[456] = 1'b0 ^~ inbuffer_data[456];
assign xnor3[457] = 1'b0 ^~ inbuffer_data[457];
assign xnor3[458] = 1'b0 ^~ inbuffer_data[458];
assign xnor3[459] = 1'b0 ^~ inbuffer_data[459];
assign xnor3[460] = 1'b0 ^~ inbuffer_data[460];
assign xnor3[461] = 1'b1 ^~ inbuffer_data[461];
assign xnor3[462] = 1'b0 ^~ inbuffer_data[462];
assign xnor3[463] = 1'b0 ^~ inbuffer_data[463];
assign xnor3[464] = 1'b0 ^~ inbuffer_data[464];
assign xnor3[465] = 1'b1 ^~ inbuffer_data[465];
assign xnor3[466] = 1'b1 ^~ inbuffer_data[466];
assign xnor3[467] = 1'b1 ^~ inbuffer_data[467];
assign xnor3[468] = 1'b1 ^~ inbuffer_data[468];
assign xnor3[469] = 1'b0 ^~ inbuffer_data[469];
assign xnor3[470] = 1'b1 ^~ inbuffer_data[470];
assign xnor3[471] = 1'b1 ^~ inbuffer_data[471];
assign xnor3[472] = 1'b1 ^~ inbuffer_data[472];
assign xnor3[473] = 1'b0 ^~ inbuffer_data[473];
assign xnor3[474] = 1'b0 ^~ inbuffer_data[474];
assign xnor3[475] = 1'b1 ^~ inbuffer_data[475];
assign xnor3[476] = 1'b1 ^~ inbuffer_data[476];
assign xnor3[477] = 1'b1 ^~ inbuffer_data[477];
assign xnor3[478] = 1'b1 ^~ inbuffer_data[478];
assign xnor3[479] = 1'b1 ^~ inbuffer_data[479];
assign xnor3[480] = 1'b1 ^~ inbuffer_data[480];
assign xnor3[481] = 1'b1 ^~ inbuffer_data[481];
assign xnor3[482] = 1'b0 ^~ inbuffer_data[482];
assign xnor3[483] = 1'b0 ^~ inbuffer_data[483];
assign xnor3[484] = 1'b0 ^~ inbuffer_data[484];
assign xnor3[485] = 1'b0 ^~ inbuffer_data[485];
assign xnor3[486] = 1'b0 ^~ inbuffer_data[486];
assign xnor3[487] = 1'b0 ^~ inbuffer_data[487];
assign xnor3[488] = 1'b0 ^~ inbuffer_data[488];
assign xnor3[489] = 1'b0 ^~ inbuffer_data[489];
assign xnor3[490] = 1'b0 ^~ inbuffer_data[490];
assign xnor3[491] = 1'b0 ^~ inbuffer_data[491];
assign xnor3[492] = 1'b0 ^~ inbuffer_data[492];
assign xnor3[493] = 1'b1 ^~ inbuffer_data[493];
assign xnor3[494] = 1'b1 ^~ inbuffer_data[494];
assign xnor3[495] = 1'b1 ^~ inbuffer_data[495];
assign xnor3[496] = 1'b0 ^~ inbuffer_data[496];
assign xnor3[497] = 1'b0 ^~ inbuffer_data[497];
assign xnor3[498] = 1'b1 ^~ inbuffer_data[498];
assign xnor3[499] = 1'b1 ^~ inbuffer_data[499];
assign xnor3[500] = 1'b0 ^~ inbuffer_data[500];
assign xnor3[501] = 1'b0 ^~ inbuffer_data[501];
assign xnor3[502] = 1'b1 ^~ inbuffer_data[502];
assign xnor3[503] = 1'b1 ^~ inbuffer_data[503];
assign xnor3[504] = 1'b1 ^~ inbuffer_data[504];
assign xnor3[505] = 1'b0 ^~ inbuffer_data[505];
assign xnor3[506] = 1'b0 ^~ inbuffer_data[506];
assign xnor3[507] = 1'b1 ^~ inbuffer_data[507];
assign xnor3[508] = 1'b1 ^~ inbuffer_data[508];
assign xnor3[509] = 1'b1 ^~ inbuffer_data[509];
assign xnor3[510] = 1'b1 ^~ inbuffer_data[510];
assign xnor3[511] = 1'b0 ^~ inbuffer_data[511];
assign xnor3[512] = 1'b0 ^~ inbuffer_data[512];
assign xnor3[513] = 1'b0 ^~ inbuffer_data[513];
assign xnor3[514] = 1'b0 ^~ inbuffer_data[514];
assign xnor3[515] = 1'b0 ^~ inbuffer_data[515];
assign xnor3[516] = 1'b0 ^~ inbuffer_data[516];
assign xnor3[517] = 1'b0 ^~ inbuffer_data[517];
assign xnor3[518] = 1'b0 ^~ inbuffer_data[518];
assign xnor3[519] = 1'b1 ^~ inbuffer_data[519];
assign xnor3[520] = 1'b1 ^~ inbuffer_data[520];
assign xnor3[521] = 1'b1 ^~ inbuffer_data[521];
assign xnor3[522] = 1'b1 ^~ inbuffer_data[522];
assign xnor3[523] = 1'b1 ^~ inbuffer_data[523];
assign xnor3[524] = 1'b0 ^~ inbuffer_data[524];
assign xnor3[525] = 1'b1 ^~ inbuffer_data[525];
assign xnor3[526] = 1'b1 ^~ inbuffer_data[526];
assign xnor3[527] = 1'b1 ^~ inbuffer_data[527];
assign xnor3[528] = 1'b0 ^~ inbuffer_data[528];
assign xnor3[529] = 1'b0 ^~ inbuffer_data[529];
assign xnor3[530] = 1'b0 ^~ inbuffer_data[530];
assign xnor3[531] = 1'b0 ^~ inbuffer_data[531];
assign xnor3[532] = 1'b1 ^~ inbuffer_data[532];
assign xnor3[533] = 1'b0 ^~ inbuffer_data[533];
assign xnor3[534] = 1'b0 ^~ inbuffer_data[534];
assign xnor3[535] = 1'b1 ^~ inbuffer_data[535];
assign xnor3[536] = 1'b1 ^~ inbuffer_data[536];
assign xnor3[537] = 1'b1 ^~ inbuffer_data[537];
assign xnor3[538] = 1'b1 ^~ inbuffer_data[538];
assign xnor3[539] = 1'b0 ^~ inbuffer_data[539];
assign xnor3[540] = 1'b0 ^~ inbuffer_data[540];
assign xnor3[541] = 1'b0 ^~ inbuffer_data[541];
assign xnor3[542] = 1'b0 ^~ inbuffer_data[542];
assign xnor3[543] = 1'b0 ^~ inbuffer_data[543];
assign xnor3[544] = 1'b0 ^~ inbuffer_data[544];
assign xnor3[545] = 1'b0 ^~ inbuffer_data[545];
assign xnor3[546] = 1'b1 ^~ inbuffer_data[546];
assign xnor3[547] = 1'b0 ^~ inbuffer_data[547];
assign xnor3[548] = 1'b1 ^~ inbuffer_data[548];
assign xnor3[549] = 1'b1 ^~ inbuffer_data[549];
assign xnor3[550] = 1'b1 ^~ inbuffer_data[550];
assign xnor3[551] = 1'b1 ^~ inbuffer_data[551];
assign xnor3[552] = 1'b1 ^~ inbuffer_data[552];
assign xnor3[553] = 1'b1 ^~ inbuffer_data[553];
assign xnor3[554] = 1'b1 ^~ inbuffer_data[554];
assign xnor3[555] = 1'b1 ^~ inbuffer_data[555];
assign xnor3[556] = 1'b0 ^~ inbuffer_data[556];
assign xnor3[557] = 1'b0 ^~ inbuffer_data[557];
assign xnor3[558] = 1'b0 ^~ inbuffer_data[558];
assign xnor3[559] = 1'b1 ^~ inbuffer_data[559];
assign xnor3[560] = 1'b0 ^~ inbuffer_data[560];
assign xnor3[561] = 1'b1 ^~ inbuffer_data[561];
assign xnor3[562] = 1'b0 ^~ inbuffer_data[562];
assign xnor3[563] = 1'b1 ^~ inbuffer_data[563];
assign xnor3[564] = 1'b1 ^~ inbuffer_data[564];
assign xnor3[565] = 1'b1 ^~ inbuffer_data[565];
assign xnor3[566] = 1'b1 ^~ inbuffer_data[566];
assign xnor3[567] = 1'b1 ^~ inbuffer_data[567];
assign xnor3[568] = 1'b1 ^~ inbuffer_data[568];
assign xnor3[569] = 1'b0 ^~ inbuffer_data[569];
assign xnor3[570] = 1'b0 ^~ inbuffer_data[570];
assign xnor3[571] = 1'b0 ^~ inbuffer_data[571];
assign xnor3[572] = 1'b0 ^~ inbuffer_data[572];
assign xnor3[573] = 1'b0 ^~ inbuffer_data[573];
assign xnor3[574] = 1'b1 ^~ inbuffer_data[574];
assign xnor3[575] = 1'b1 ^~ inbuffer_data[575];
assign xnor3[576] = 1'b1 ^~ inbuffer_data[576];
assign xnor3[577] = 1'b1 ^~ inbuffer_data[577];
assign xnor3[578] = 1'b1 ^~ inbuffer_data[578];
assign xnor3[579] = 1'b1 ^~ inbuffer_data[579];
assign xnor3[580] = 1'b1 ^~ inbuffer_data[580];
assign xnor3[581] = 1'b1 ^~ inbuffer_data[581];
assign xnor3[582] = 1'b0 ^~ inbuffer_data[582];
assign xnor3[583] = 1'b0 ^~ inbuffer_data[583];
assign xnor3[584] = 1'b0 ^~ inbuffer_data[584];
assign xnor3[585] = 1'b1 ^~ inbuffer_data[585];
assign xnor3[586] = 1'b0 ^~ inbuffer_data[586];
assign xnor3[587] = 1'b0 ^~ inbuffer_data[587];
assign xnor3[588] = 1'b0 ^~ inbuffer_data[588];
assign xnor3[589] = 1'b1 ^~ inbuffer_data[589];
assign xnor3[590] = 1'b0 ^~ inbuffer_data[590];
assign xnor3[591] = 1'b1 ^~ inbuffer_data[591];
assign xnor3[592] = 1'b1 ^~ inbuffer_data[592];
assign xnor3[593] = 1'b1 ^~ inbuffer_data[593];
assign xnor3[594] = 1'b1 ^~ inbuffer_data[594];
assign xnor3[595] = 1'b1 ^~ inbuffer_data[595];
assign xnor3[596] = 1'b1 ^~ inbuffer_data[596];
assign xnor3[597] = 1'b0 ^~ inbuffer_data[597];
assign xnor3[598] = 1'b0 ^~ inbuffer_data[598];
assign xnor3[599] = 1'b1 ^~ inbuffer_data[599];
assign xnor3[600] = 1'b0 ^~ inbuffer_data[600];
assign xnor3[601] = 1'b0 ^~ inbuffer_data[601];
assign xnor3[602] = 1'b0 ^~ inbuffer_data[602];
assign xnor3[603] = 1'b0 ^~ inbuffer_data[603];
assign xnor3[604] = 1'b0 ^~ inbuffer_data[604];
assign xnor3[605] = 1'b1 ^~ inbuffer_data[605];
assign xnor3[606] = 1'b1 ^~ inbuffer_data[606];
assign xnor3[607] = 1'b1 ^~ inbuffer_data[607];
assign xnor3[608] = 1'b0 ^~ inbuffer_data[608];
assign xnor3[609] = 1'b1 ^~ inbuffer_data[609];
assign xnor3[610] = 1'b1 ^~ inbuffer_data[610];
assign xnor3[611] = 1'b0 ^~ inbuffer_data[611];
assign xnor3[612] = 1'b0 ^~ inbuffer_data[612];
assign xnor3[613] = 1'b0 ^~ inbuffer_data[613];
assign xnor3[614] = 1'b0 ^~ inbuffer_data[614];
assign xnor3[615] = 1'b0 ^~ inbuffer_data[615];
assign xnor3[616] = 1'b0 ^~ inbuffer_data[616];
assign xnor3[617] = 1'b0 ^~ inbuffer_data[617];
assign xnor3[618] = 1'b1 ^~ inbuffer_data[618];
assign xnor3[619] = 1'b1 ^~ inbuffer_data[619];
assign xnor3[620] = 1'b1 ^~ inbuffer_data[620];
assign xnor3[621] = 1'b0 ^~ inbuffer_data[621];
assign xnor3[622] = 1'b1 ^~ inbuffer_data[622];
assign xnor3[623] = 1'b1 ^~ inbuffer_data[623];
assign xnor3[624] = 1'b0 ^~ inbuffer_data[624];
assign xnor3[625] = 1'b1 ^~ inbuffer_data[625];
assign xnor3[626] = 1'b0 ^~ inbuffer_data[626];
assign xnor3[627] = 1'b1 ^~ inbuffer_data[627];
assign xnor3[628] = 1'b1 ^~ inbuffer_data[628];
assign xnor3[629] = 1'b0 ^~ inbuffer_data[629];
assign xnor3[630] = 1'b1 ^~ inbuffer_data[630];
assign xnor3[631] = 1'b0 ^~ inbuffer_data[631];
assign xnor3[632] = 1'b1 ^~ inbuffer_data[632];
assign xnor3[633] = 1'b1 ^~ inbuffer_data[633];
assign xnor3[634] = 1'b1 ^~ inbuffer_data[634];
assign xnor3[635] = 1'b1 ^~ inbuffer_data[635];
assign xnor3[636] = 1'b1 ^~ inbuffer_data[636];
assign xnor3[637] = 1'b0 ^~ inbuffer_data[637];
assign xnor3[638] = 1'b0 ^~ inbuffer_data[638];
assign xnor3[639] = 1'b0 ^~ inbuffer_data[639];
assign xnor3[640] = 1'b1 ^~ inbuffer_data[640];
assign xnor3[641] = 1'b0 ^~ inbuffer_data[641];
assign xnor3[642] = 1'b1 ^~ inbuffer_data[642];
assign xnor3[643] = 1'b1 ^~ inbuffer_data[643];
assign xnor3[644] = 1'b0 ^~ inbuffer_data[644];
assign xnor3[645] = 1'b0 ^~ inbuffer_data[645];
assign xnor3[646] = 1'b0 ^~ inbuffer_data[646];
assign xnor3[647] = 1'b1 ^~ inbuffer_data[647];
assign xnor3[648] = 1'b1 ^~ inbuffer_data[648];
assign xnor3[649] = 1'b1 ^~ inbuffer_data[649];
assign xnor3[650] = 1'b1 ^~ inbuffer_data[650];
assign xnor3[651] = 1'b1 ^~ inbuffer_data[651];
assign xnor3[652] = 1'b1 ^~ inbuffer_data[652];
assign xnor3[653] = 1'b1 ^~ inbuffer_data[653];
assign xnor3[654] = 1'b1 ^~ inbuffer_data[654];
assign xnor3[655] = 1'b1 ^~ inbuffer_data[655];
assign xnor3[656] = 1'b0 ^~ inbuffer_data[656];
assign xnor3[657] = 1'b0 ^~ inbuffer_data[657];
assign xnor3[658] = 1'b0 ^~ inbuffer_data[658];
assign xnor3[659] = 1'b0 ^~ inbuffer_data[659];
assign xnor3[660] = 1'b0 ^~ inbuffer_data[660];
assign xnor3[661] = 1'b1 ^~ inbuffer_data[661];
assign xnor3[662] = 1'b1 ^~ inbuffer_data[662];
assign xnor3[663] = 1'b0 ^~ inbuffer_data[663];
assign xnor3[664] = 1'b1 ^~ inbuffer_data[664];
assign xnor3[665] = 1'b0 ^~ inbuffer_data[665];
assign xnor3[666] = 1'b0 ^~ inbuffer_data[666];
assign xnor3[667] = 1'b0 ^~ inbuffer_data[667];
assign xnor3[668] = 1'b1 ^~ inbuffer_data[668];
assign xnor3[669] = 1'b0 ^~ inbuffer_data[669];
assign xnor3[670] = 1'b0 ^~ inbuffer_data[670];
assign xnor3[671] = 1'b0 ^~ inbuffer_data[671];
assign xnor3[672] = 1'b1 ^~ inbuffer_data[672];
assign xnor3[673] = 1'b0 ^~ inbuffer_data[673];
assign xnor3[674] = 1'b0 ^~ inbuffer_data[674];
assign xnor3[675] = 1'b1 ^~ inbuffer_data[675];
assign xnor3[676] = 1'b1 ^~ inbuffer_data[676];
assign xnor3[677] = 1'b1 ^~ inbuffer_data[677];
assign xnor3[678] = 1'b1 ^~ inbuffer_data[678];
assign xnor3[679] = 1'b1 ^~ inbuffer_data[679];
assign xnor3[680] = 1'b1 ^~ inbuffer_data[680];
assign xnor3[681] = 1'b1 ^~ inbuffer_data[681];
assign xnor3[682] = 1'b1 ^~ inbuffer_data[682];
assign xnor3[683] = 1'b1 ^~ inbuffer_data[683];
assign xnor3[684] = 1'b1 ^~ inbuffer_data[684];
assign xnor3[685] = 1'b1 ^~ inbuffer_data[685];
assign xnor3[686] = 1'b1 ^~ inbuffer_data[686];
assign xnor3[687] = 1'b0 ^~ inbuffer_data[687];
assign xnor3[688] = 1'b1 ^~ inbuffer_data[688];
assign xnor3[689] = 1'b1 ^~ inbuffer_data[689];
assign xnor3[690] = 1'b0 ^~ inbuffer_data[690];
assign xnor3[691] = 1'b0 ^~ inbuffer_data[691];
assign xnor3[692] = 1'b0 ^~ inbuffer_data[692];
assign xnor3[693] = 1'b1 ^~ inbuffer_data[693];
assign xnor3[694] = 1'b0 ^~ inbuffer_data[694];
assign xnor3[695] = 1'b1 ^~ inbuffer_data[695];
assign xnor3[696] = 1'b0 ^~ inbuffer_data[696];
assign xnor3[697] = 1'b1 ^~ inbuffer_data[697];
assign xnor3[698] = 1'b1 ^~ inbuffer_data[698];
assign xnor3[699] = 1'b0 ^~ inbuffer_data[699];
assign xnor3[700] = 1'b1 ^~ inbuffer_data[700];
assign xnor3[701] = 1'b0 ^~ inbuffer_data[701];
assign xnor3[702] = 1'b0 ^~ inbuffer_data[702];
assign xnor3[703] = 1'b1 ^~ inbuffer_data[703];
assign xnor3[704] = 1'b0 ^~ inbuffer_data[704];
assign xnor3[705] = 1'b0 ^~ inbuffer_data[705];
assign xnor3[706] = 1'b1 ^~ inbuffer_data[706];
assign xnor3[707] = 1'b1 ^~ inbuffer_data[707];
assign xnor3[708] = 1'b1 ^~ inbuffer_data[708];
assign xnor3[709] = 1'b1 ^~ inbuffer_data[709];
assign xnor3[710] = 1'b1 ^~ inbuffer_data[710];
assign xnor3[711] = 1'b1 ^~ inbuffer_data[711];
assign xnor3[712] = 1'b1 ^~ inbuffer_data[712];
assign xnor3[713] = 1'b1 ^~ inbuffer_data[713];
assign xnor3[714] = 1'b1 ^~ inbuffer_data[714];
assign xnor3[715] = 1'b1 ^~ inbuffer_data[715];
assign xnor3[716] = 1'b1 ^~ inbuffer_data[716];
assign xnor3[717] = 1'b1 ^~ inbuffer_data[717];
assign xnor3[718] = 1'b1 ^~ inbuffer_data[718];
assign xnor3[719] = 1'b0 ^~ inbuffer_data[719];
assign xnor3[720] = 1'b1 ^~ inbuffer_data[720];
assign xnor3[721] = 1'b0 ^~ inbuffer_data[721];
assign xnor3[722] = 1'b0 ^~ inbuffer_data[722];
assign xnor3[723] = 1'b0 ^~ inbuffer_data[723];
assign xnor3[724] = 1'b1 ^~ inbuffer_data[724];
assign xnor3[725] = 1'b0 ^~ inbuffer_data[725];
assign xnor3[726] = 1'b0 ^~ inbuffer_data[726];
assign xnor3[727] = 1'b0 ^~ inbuffer_data[727];
assign xnor3[728] = 1'b0 ^~ inbuffer_data[728];
assign xnor3[729] = 1'b0 ^~ inbuffer_data[729];
assign xnor3[730] = 1'b1 ^~ inbuffer_data[730];
assign xnor3[731] = 1'b1 ^~ inbuffer_data[731];
assign xnor3[732] = 1'b0 ^~ inbuffer_data[732];
assign xnor3[733] = 1'b1 ^~ inbuffer_data[733];
assign xnor3[734] = 1'b0 ^~ inbuffer_data[734];
assign xnor3[735] = 1'b1 ^~ inbuffer_data[735];
assign xnor3[736] = 1'b0 ^~ inbuffer_data[736];
assign xnor3[737] = 1'b0 ^~ inbuffer_data[737];
assign xnor3[738] = 1'b0 ^~ inbuffer_data[738];
assign xnor3[739] = 1'b0 ^~ inbuffer_data[739];
assign xnor3[740] = 1'b0 ^~ inbuffer_data[740];
assign xnor3[741] = 1'b0 ^~ inbuffer_data[741];
assign xnor3[742] = 1'b1 ^~ inbuffer_data[742];
assign xnor3[743] = 1'b0 ^~ inbuffer_data[743];
assign xnor3[744] = 1'b1 ^~ inbuffer_data[744];
assign xnor3[745] = 1'b0 ^~ inbuffer_data[745];
assign xnor3[746] = 1'b1 ^~ inbuffer_data[746];
assign xnor3[747] = 1'b1 ^~ inbuffer_data[747];
assign xnor3[748] = 1'b1 ^~ inbuffer_data[748];
assign xnor3[749] = 1'b0 ^~ inbuffer_data[749];
assign xnor3[750] = 1'b0 ^~ inbuffer_data[750];
assign xnor3[751] = 1'b0 ^~ inbuffer_data[751];
assign xnor3[752] = 1'b1 ^~ inbuffer_data[752];
assign xnor3[753] = 1'b1 ^~ inbuffer_data[753];
assign xnor3[754] = 1'b1 ^~ inbuffer_data[754];
assign xnor3[755] = 1'b0 ^~ inbuffer_data[755];
assign xnor3[756] = 1'b0 ^~ inbuffer_data[756];
assign xnor3[757] = 1'b0 ^~ inbuffer_data[757];
assign xnor3[758] = 1'b1 ^~ inbuffer_data[758];
assign xnor3[759] = 1'b1 ^~ inbuffer_data[759];
assign xnor3[760] = 1'b1 ^~ inbuffer_data[760];
assign xnor3[761] = 1'b0 ^~ inbuffer_data[761];
assign xnor3[762] = 1'b1 ^~ inbuffer_data[762];
assign xnor3[763] = 1'b0 ^~ inbuffer_data[763];
assign xnor3[764] = 1'b1 ^~ inbuffer_data[764];
assign xnor3[765] = 1'b0 ^~ inbuffer_data[765];
assign xnor3[766] = 1'b1 ^~ inbuffer_data[766];
assign xnor3[767] = 1'b1 ^~ inbuffer_data[767];
assign xnor3[768] = 1'b0 ^~ inbuffer_data[768];
assign xnor3[769] = 1'b0 ^~ inbuffer_data[769];
assign xnor3[770] = 1'b0 ^~ inbuffer_data[770];
assign xnor3[771] = 1'b0 ^~ inbuffer_data[771];
assign xnor3[772] = 1'b0 ^~ inbuffer_data[772];
assign xnor3[773] = 1'b1 ^~ inbuffer_data[773];
assign xnor3[774] = 1'b1 ^~ inbuffer_data[774];
assign xnor3[775] = 1'b1 ^~ inbuffer_data[775];
assign xnor3[776] = 1'b1 ^~ inbuffer_data[776];
assign xnor3[777] = 1'b0 ^~ inbuffer_data[777];
assign xnor3[778] = 1'b1 ^~ inbuffer_data[778];
assign xnor3[779] = 1'b1 ^~ inbuffer_data[779];
assign xnor3[780] = 1'b0 ^~ inbuffer_data[780];
assign xnor3[781] = 1'b1 ^~ inbuffer_data[781];
assign xnor3[782] = 1'b0 ^~ inbuffer_data[782];
assign xnor3[783] = 1'b1 ^~ inbuffer_data[783];
assign xnor4[0] = 1'b1 ^~ inbuffer_data[0];
assign xnor4[1] = 1'b1 ^~ inbuffer_data[1];
assign xnor4[2] = 1'b0 ^~ inbuffer_data[2];
assign xnor4[3] = 1'b1 ^~ inbuffer_data[3];
assign xnor4[4] = 1'b1 ^~ inbuffer_data[4];
assign xnor4[5] = 1'b1 ^~ inbuffer_data[5];
assign xnor4[6] = 1'b1 ^~ inbuffer_data[6];
assign xnor4[7] = 1'b1 ^~ inbuffer_data[7];
assign xnor4[8] = 1'b0 ^~ inbuffer_data[8];
assign xnor4[9] = 1'b1 ^~ inbuffer_data[9];
assign xnor4[10] = 1'b0 ^~ inbuffer_data[10];
assign xnor4[11] = 1'b1 ^~ inbuffer_data[11];
assign xnor4[12] = 1'b0 ^~ inbuffer_data[12];
assign xnor4[13] = 1'b0 ^~ inbuffer_data[13];
assign xnor4[14] = 1'b1 ^~ inbuffer_data[14];
assign xnor4[15] = 1'b0 ^~ inbuffer_data[15];
assign xnor4[16] = 1'b1 ^~ inbuffer_data[16];
assign xnor4[17] = 1'b0 ^~ inbuffer_data[17];
assign xnor4[18] = 1'b0 ^~ inbuffer_data[18];
assign xnor4[19] = 1'b0 ^~ inbuffer_data[19];
assign xnor4[20] = 1'b0 ^~ inbuffer_data[20];
assign xnor4[21] = 1'b1 ^~ inbuffer_data[21];
assign xnor4[22] = 1'b1 ^~ inbuffer_data[22];
assign xnor4[23] = 1'b0 ^~ inbuffer_data[23];
assign xnor4[24] = 1'b1 ^~ inbuffer_data[24];
assign xnor4[25] = 1'b1 ^~ inbuffer_data[25];
assign xnor4[26] = 1'b1 ^~ inbuffer_data[26];
assign xnor4[27] = 1'b0 ^~ inbuffer_data[27];
assign xnor4[28] = 1'b0 ^~ inbuffer_data[28];
assign xnor4[29] = 1'b1 ^~ inbuffer_data[29];
assign xnor4[30] = 1'b1 ^~ inbuffer_data[30];
assign xnor4[31] = 1'b0 ^~ inbuffer_data[31];
assign xnor4[32] = 1'b1 ^~ inbuffer_data[32];
assign xnor4[33] = 1'b1 ^~ inbuffer_data[33];
assign xnor4[34] = 1'b1 ^~ inbuffer_data[34];
assign xnor4[35] = 1'b0 ^~ inbuffer_data[35];
assign xnor4[36] = 1'b0 ^~ inbuffer_data[36];
assign xnor4[37] = 1'b0 ^~ inbuffer_data[37];
assign xnor4[38] = 1'b0 ^~ inbuffer_data[38];
assign xnor4[39] = 1'b0 ^~ inbuffer_data[39];
assign xnor4[40] = 1'b1 ^~ inbuffer_data[40];
assign xnor4[41] = 1'b1 ^~ inbuffer_data[41];
assign xnor4[42] = 1'b0 ^~ inbuffer_data[42];
assign xnor4[43] = 1'b0 ^~ inbuffer_data[43];
assign xnor4[44] = 1'b1 ^~ inbuffer_data[44];
assign xnor4[45] = 1'b1 ^~ inbuffer_data[45];
assign xnor4[46] = 1'b0 ^~ inbuffer_data[46];
assign xnor4[47] = 1'b1 ^~ inbuffer_data[47];
assign xnor4[48] = 1'b1 ^~ inbuffer_data[48];
assign xnor4[49] = 1'b0 ^~ inbuffer_data[49];
assign xnor4[50] = 1'b1 ^~ inbuffer_data[50];
assign xnor4[51] = 1'b0 ^~ inbuffer_data[51];
assign xnor4[52] = 1'b1 ^~ inbuffer_data[52];
assign xnor4[53] = 1'b1 ^~ inbuffer_data[53];
assign xnor4[54] = 1'b0 ^~ inbuffer_data[54];
assign xnor4[55] = 1'b1 ^~ inbuffer_data[55];
assign xnor4[56] = 1'b1 ^~ inbuffer_data[56];
assign xnor4[57] = 1'b0 ^~ inbuffer_data[57];
assign xnor4[58] = 1'b0 ^~ inbuffer_data[58];
assign xnor4[59] = 1'b0 ^~ inbuffer_data[59];
assign xnor4[60] = 1'b0 ^~ inbuffer_data[60];
assign xnor4[61] = 1'b1 ^~ inbuffer_data[61];
assign xnor4[62] = 1'b0 ^~ inbuffer_data[62];
assign xnor4[63] = 1'b1 ^~ inbuffer_data[63];
assign xnor4[64] = 1'b0 ^~ inbuffer_data[64];
assign xnor4[65] = 1'b0 ^~ inbuffer_data[65];
assign xnor4[66] = 1'b0 ^~ inbuffer_data[66];
assign xnor4[67] = 1'b0 ^~ inbuffer_data[67];
assign xnor4[68] = 1'b1 ^~ inbuffer_data[68];
assign xnor4[69] = 1'b1 ^~ inbuffer_data[69];
assign xnor4[70] = 1'b0 ^~ inbuffer_data[70];
assign xnor4[71] = 1'b0 ^~ inbuffer_data[71];
assign xnor4[72] = 1'b0 ^~ inbuffer_data[72];
assign xnor4[73] = 1'b0 ^~ inbuffer_data[73];
assign xnor4[74] = 1'b0 ^~ inbuffer_data[74];
assign xnor4[75] = 1'b0 ^~ inbuffer_data[75];
assign xnor4[76] = 1'b1 ^~ inbuffer_data[76];
assign xnor4[77] = 1'b1 ^~ inbuffer_data[77];
assign xnor4[78] = 1'b1 ^~ inbuffer_data[78];
assign xnor4[79] = 1'b1 ^~ inbuffer_data[79];
assign xnor4[80] = 1'b0 ^~ inbuffer_data[80];
assign xnor4[81] = 1'b1 ^~ inbuffer_data[81];
assign xnor4[82] = 1'b1 ^~ inbuffer_data[82];
assign xnor4[83] = 1'b1 ^~ inbuffer_data[83];
assign xnor4[84] = 1'b1 ^~ inbuffer_data[84];
assign xnor4[85] = 1'b1 ^~ inbuffer_data[85];
assign xnor4[86] = 1'b1 ^~ inbuffer_data[86];
assign xnor4[87] = 1'b1 ^~ inbuffer_data[87];
assign xnor4[88] = 1'b1 ^~ inbuffer_data[88];
assign xnor4[89] = 1'b1 ^~ inbuffer_data[89];
assign xnor4[90] = 1'b0 ^~ inbuffer_data[90];
assign xnor4[91] = 1'b0 ^~ inbuffer_data[91];
assign xnor4[92] = 1'b0 ^~ inbuffer_data[92];
assign xnor4[93] = 1'b0 ^~ inbuffer_data[93];
assign xnor4[94] = 1'b0 ^~ inbuffer_data[94];
assign xnor4[95] = 1'b0 ^~ inbuffer_data[95];
assign xnor4[96] = 1'b0 ^~ inbuffer_data[96];
assign xnor4[97] = 1'b0 ^~ inbuffer_data[97];
assign xnor4[98] = 1'b0 ^~ inbuffer_data[98];
assign xnor4[99] = 1'b0 ^~ inbuffer_data[99];
assign xnor4[100] = 1'b0 ^~ inbuffer_data[100];
assign xnor4[101] = 1'b0 ^~ inbuffer_data[101];
assign xnor4[102] = 1'b0 ^~ inbuffer_data[102];
assign xnor4[103] = 1'b0 ^~ inbuffer_data[103];
assign xnor4[104] = 1'b1 ^~ inbuffer_data[104];
assign xnor4[105] = 1'b0 ^~ inbuffer_data[105];
assign xnor4[106] = 1'b1 ^~ inbuffer_data[106];
assign xnor4[107] = 1'b1 ^~ inbuffer_data[107];
assign xnor4[108] = 1'b0 ^~ inbuffer_data[108];
assign xnor4[109] = 1'b1 ^~ inbuffer_data[109];
assign xnor4[110] = 1'b1 ^~ inbuffer_data[110];
assign xnor4[111] = 1'b1 ^~ inbuffer_data[111];
assign xnor4[112] = 1'b0 ^~ inbuffer_data[112];
assign xnor4[113] = 1'b1 ^~ inbuffer_data[113];
assign xnor4[114] = 1'b1 ^~ inbuffer_data[114];
assign xnor4[115] = 1'b1 ^~ inbuffer_data[115];
assign xnor4[116] = 1'b1 ^~ inbuffer_data[116];
assign xnor4[117] = 1'b1 ^~ inbuffer_data[117];
assign xnor4[118] = 1'b0 ^~ inbuffer_data[118];
assign xnor4[119] = 1'b0 ^~ inbuffer_data[119];
assign xnor4[120] = 1'b1 ^~ inbuffer_data[120];
assign xnor4[121] = 1'b0 ^~ inbuffer_data[121];
assign xnor4[122] = 1'b0 ^~ inbuffer_data[122];
assign xnor4[123] = 1'b0 ^~ inbuffer_data[123];
assign xnor4[124] = 1'b0 ^~ inbuffer_data[124];
assign xnor4[125] = 1'b0 ^~ inbuffer_data[125];
assign xnor4[126] = 1'b0 ^~ inbuffer_data[126];
assign xnor4[127] = 1'b0 ^~ inbuffer_data[127];
assign xnor4[128] = 1'b0 ^~ inbuffer_data[128];
assign xnor4[129] = 1'b1 ^~ inbuffer_data[129];
assign xnor4[130] = 1'b0 ^~ inbuffer_data[130];
assign xnor4[131] = 1'b1 ^~ inbuffer_data[131];
assign xnor4[132] = 1'b1 ^~ inbuffer_data[132];
assign xnor4[133] = 1'b1 ^~ inbuffer_data[133];
assign xnor4[134] = 1'b1 ^~ inbuffer_data[134];
assign xnor4[135] = 1'b1 ^~ inbuffer_data[135];
assign xnor4[136] = 1'b1 ^~ inbuffer_data[136];
assign xnor4[137] = 1'b1 ^~ inbuffer_data[137];
assign xnor4[138] = 1'b0 ^~ inbuffer_data[138];
assign xnor4[139] = 1'b1 ^~ inbuffer_data[139];
assign xnor4[140] = 1'b0 ^~ inbuffer_data[140];
assign xnor4[141] = 1'b1 ^~ inbuffer_data[141];
assign xnor4[142] = 1'b1 ^~ inbuffer_data[142];
assign xnor4[143] = 1'b0 ^~ inbuffer_data[143];
assign xnor4[144] = 1'b0 ^~ inbuffer_data[144];
assign xnor4[145] = 1'b1 ^~ inbuffer_data[145];
assign xnor4[146] = 1'b0 ^~ inbuffer_data[146];
assign xnor4[147] = 1'b1 ^~ inbuffer_data[147];
assign xnor4[148] = 1'b1 ^~ inbuffer_data[148];
assign xnor4[149] = 1'b1 ^~ inbuffer_data[149];
assign xnor4[150] = 1'b0 ^~ inbuffer_data[150];
assign xnor4[151] = 1'b0 ^~ inbuffer_data[151];
assign xnor4[152] = 1'b1 ^~ inbuffer_data[152];
assign xnor4[153] = 1'b0 ^~ inbuffer_data[153];
assign xnor4[154] = 1'b1 ^~ inbuffer_data[154];
assign xnor4[155] = 1'b0 ^~ inbuffer_data[155];
assign xnor4[156] = 1'b0 ^~ inbuffer_data[156];
assign xnor4[157] = 1'b1 ^~ inbuffer_data[157];
assign xnor4[158] = 1'b1 ^~ inbuffer_data[158];
assign xnor4[159] = 1'b1 ^~ inbuffer_data[159];
assign xnor4[160] = 1'b1 ^~ inbuffer_data[160];
assign xnor4[161] = 1'b1 ^~ inbuffer_data[161];
assign xnor4[162] = 1'b1 ^~ inbuffer_data[162];
assign xnor4[163] = 1'b1 ^~ inbuffer_data[163];
assign xnor4[164] = 1'b1 ^~ inbuffer_data[164];
assign xnor4[165] = 1'b1 ^~ inbuffer_data[165];
assign xnor4[166] = 1'b1 ^~ inbuffer_data[166];
assign xnor4[167] = 1'b0 ^~ inbuffer_data[167];
assign xnor4[168] = 1'b1 ^~ inbuffer_data[168];
assign xnor4[169] = 1'b0 ^~ inbuffer_data[169];
assign xnor4[170] = 1'b0 ^~ inbuffer_data[170];
assign xnor4[171] = 1'b1 ^~ inbuffer_data[171];
assign xnor4[172] = 1'b1 ^~ inbuffer_data[172];
assign xnor4[173] = 1'b1 ^~ inbuffer_data[173];
assign xnor4[174] = 1'b1 ^~ inbuffer_data[174];
assign xnor4[175] = 1'b1 ^~ inbuffer_data[175];
assign xnor4[176] = 1'b0 ^~ inbuffer_data[176];
assign xnor4[177] = 1'b1 ^~ inbuffer_data[177];
assign xnor4[178] = 1'b1 ^~ inbuffer_data[178];
assign xnor4[179] = 1'b0 ^~ inbuffer_data[179];
assign xnor4[180] = 1'b0 ^~ inbuffer_data[180];
assign xnor4[181] = 1'b0 ^~ inbuffer_data[181];
assign xnor4[182] = 1'b0 ^~ inbuffer_data[182];
assign xnor4[183] = 1'b0 ^~ inbuffer_data[183];
assign xnor4[184] = 1'b0 ^~ inbuffer_data[184];
assign xnor4[185] = 1'b0 ^~ inbuffer_data[185];
assign xnor4[186] = 1'b0 ^~ inbuffer_data[186];
assign xnor4[187] = 1'b0 ^~ inbuffer_data[187];
assign xnor4[188] = 1'b1 ^~ inbuffer_data[188];
assign xnor4[189] = 1'b1 ^~ inbuffer_data[189];
assign xnor4[190] = 1'b1 ^~ inbuffer_data[190];
assign xnor4[191] = 1'b1 ^~ inbuffer_data[191];
assign xnor4[192] = 1'b1 ^~ inbuffer_data[192];
assign xnor4[193] = 1'b0 ^~ inbuffer_data[193];
assign xnor4[194] = 1'b1 ^~ inbuffer_data[194];
assign xnor4[195] = 1'b1 ^~ inbuffer_data[195];
assign xnor4[196] = 1'b0 ^~ inbuffer_data[196];
assign xnor4[197] = 1'b1 ^~ inbuffer_data[197];
assign xnor4[198] = 1'b1 ^~ inbuffer_data[198];
assign xnor4[199] = 1'b1 ^~ inbuffer_data[199];
assign xnor4[200] = 1'b1 ^~ inbuffer_data[200];
assign xnor4[201] = 1'b1 ^~ inbuffer_data[201];
assign xnor4[202] = 1'b0 ^~ inbuffer_data[202];
assign xnor4[203] = 1'b0 ^~ inbuffer_data[203];
assign xnor4[204] = 1'b1 ^~ inbuffer_data[204];
assign xnor4[205] = 1'b0 ^~ inbuffer_data[205];
assign xnor4[206] = 1'b1 ^~ inbuffer_data[206];
assign xnor4[207] = 1'b0 ^~ inbuffer_data[207];
assign xnor4[208] = 1'b0 ^~ inbuffer_data[208];
assign xnor4[209] = 1'b0 ^~ inbuffer_data[209];
assign xnor4[210] = 1'b0 ^~ inbuffer_data[210];
assign xnor4[211] = 1'b0 ^~ inbuffer_data[211];
assign xnor4[212] = 1'b0 ^~ inbuffer_data[212];
assign xnor4[213] = 1'b0 ^~ inbuffer_data[213];
assign xnor4[214] = 1'b1 ^~ inbuffer_data[214];
assign xnor4[215] = 1'b0 ^~ inbuffer_data[215];
assign xnor4[216] = 1'b1 ^~ inbuffer_data[216];
assign xnor4[217] = 1'b1 ^~ inbuffer_data[217];
assign xnor4[218] = 1'b1 ^~ inbuffer_data[218];
assign xnor4[219] = 1'b1 ^~ inbuffer_data[219];
assign xnor4[220] = 1'b0 ^~ inbuffer_data[220];
assign xnor4[221] = 1'b1 ^~ inbuffer_data[221];
assign xnor4[222] = 1'b0 ^~ inbuffer_data[222];
assign xnor4[223] = 1'b1 ^~ inbuffer_data[223];
assign xnor4[224] = 1'b0 ^~ inbuffer_data[224];
assign xnor4[225] = 1'b0 ^~ inbuffer_data[225];
assign xnor4[226] = 1'b0 ^~ inbuffer_data[226];
assign xnor4[227] = 1'b1 ^~ inbuffer_data[227];
assign xnor4[228] = 1'b0 ^~ inbuffer_data[228];
assign xnor4[229] = 1'b1 ^~ inbuffer_data[229];
assign xnor4[230] = 1'b1 ^~ inbuffer_data[230];
assign xnor4[231] = 1'b0 ^~ inbuffer_data[231];
assign xnor4[232] = 1'b0 ^~ inbuffer_data[232];
assign xnor4[233] = 1'b1 ^~ inbuffer_data[233];
assign xnor4[234] = 1'b0 ^~ inbuffer_data[234];
assign xnor4[235] = 1'b0 ^~ inbuffer_data[235];
assign xnor4[236] = 1'b0 ^~ inbuffer_data[236];
assign xnor4[237] = 1'b0 ^~ inbuffer_data[237];
assign xnor4[238] = 1'b0 ^~ inbuffer_data[238];
assign xnor4[239] = 1'b0 ^~ inbuffer_data[239];
assign xnor4[240] = 1'b0 ^~ inbuffer_data[240];
assign xnor4[241] = 1'b0 ^~ inbuffer_data[241];
assign xnor4[242] = 1'b1 ^~ inbuffer_data[242];
assign xnor4[243] = 1'b1 ^~ inbuffer_data[243];
assign xnor4[244] = 1'b0 ^~ inbuffer_data[244];
assign xnor4[245] = 1'b0 ^~ inbuffer_data[245];
assign xnor4[246] = 1'b1 ^~ inbuffer_data[246];
assign xnor4[247] = 1'b1 ^~ inbuffer_data[247];
assign xnor4[248] = 1'b1 ^~ inbuffer_data[248];
assign xnor4[249] = 1'b1 ^~ inbuffer_data[249];
assign xnor4[250] = 1'b0 ^~ inbuffer_data[250];
assign xnor4[251] = 1'b0 ^~ inbuffer_data[251];
assign xnor4[252] = 1'b0 ^~ inbuffer_data[252];
assign xnor4[253] = 1'b1 ^~ inbuffer_data[253];
assign xnor4[254] = 1'b1 ^~ inbuffer_data[254];
assign xnor4[255] = 1'b0 ^~ inbuffer_data[255];
assign xnor4[256] = 1'b0 ^~ inbuffer_data[256];
assign xnor4[257] = 1'b1 ^~ inbuffer_data[257];
assign xnor4[258] = 1'b0 ^~ inbuffer_data[258];
assign xnor4[259] = 1'b1 ^~ inbuffer_data[259];
assign xnor4[260] = 1'b0 ^~ inbuffer_data[260];
assign xnor4[261] = 1'b0 ^~ inbuffer_data[261];
assign xnor4[262] = 1'b0 ^~ inbuffer_data[262];
assign xnor4[263] = 1'b0 ^~ inbuffer_data[263];
assign xnor4[264] = 1'b0 ^~ inbuffer_data[264];
assign xnor4[265] = 1'b0 ^~ inbuffer_data[265];
assign xnor4[266] = 1'b0 ^~ inbuffer_data[266];
assign xnor4[267] = 1'b0 ^~ inbuffer_data[267];
assign xnor4[268] = 1'b0 ^~ inbuffer_data[268];
assign xnor4[269] = 1'b0 ^~ inbuffer_data[269];
assign xnor4[270] = 1'b1 ^~ inbuffer_data[270];
assign xnor4[271] = 1'b0 ^~ inbuffer_data[271];
assign xnor4[272] = 1'b1 ^~ inbuffer_data[272];
assign xnor4[273] = 1'b1 ^~ inbuffer_data[273];
assign xnor4[274] = 1'b0 ^~ inbuffer_data[274];
assign xnor4[275] = 1'b0 ^~ inbuffer_data[275];
assign xnor4[276] = 1'b0 ^~ inbuffer_data[276];
assign xnor4[277] = 1'b0 ^~ inbuffer_data[277];
assign xnor4[278] = 1'b1 ^~ inbuffer_data[278];
assign xnor4[279] = 1'b0 ^~ inbuffer_data[279];
assign xnor4[280] = 1'b1 ^~ inbuffer_data[280];
assign xnor4[281] = 1'b1 ^~ inbuffer_data[281];
assign xnor4[282] = 1'b0 ^~ inbuffer_data[282];
assign xnor4[283] = 1'b1 ^~ inbuffer_data[283];
assign xnor4[284] = 1'b0 ^~ inbuffer_data[284];
assign xnor4[285] = 1'b0 ^~ inbuffer_data[285];
assign xnor4[286] = 1'b0 ^~ inbuffer_data[286];
assign xnor4[287] = 1'b0 ^~ inbuffer_data[287];
assign xnor4[288] = 1'b1 ^~ inbuffer_data[288];
assign xnor4[289] = 1'b1 ^~ inbuffer_data[289];
assign xnor4[290] = 1'b1 ^~ inbuffer_data[290];
assign xnor4[291] = 1'b1 ^~ inbuffer_data[291];
assign xnor4[292] = 1'b1 ^~ inbuffer_data[292];
assign xnor4[293] = 1'b0 ^~ inbuffer_data[293];
assign xnor4[294] = 1'b0 ^~ inbuffer_data[294];
assign xnor4[295] = 1'b0 ^~ inbuffer_data[295];
assign xnor4[296] = 1'b0 ^~ inbuffer_data[296];
assign xnor4[297] = 1'b1 ^~ inbuffer_data[297];
assign xnor4[298] = 1'b1 ^~ inbuffer_data[298];
assign xnor4[299] = 1'b1 ^~ inbuffer_data[299];
assign xnor4[300] = 1'b0 ^~ inbuffer_data[300];
assign xnor4[301] = 1'b0 ^~ inbuffer_data[301];
assign xnor4[302] = 1'b0 ^~ inbuffer_data[302];
assign xnor4[303] = 1'b0 ^~ inbuffer_data[303];
assign xnor4[304] = 1'b0 ^~ inbuffer_data[304];
assign xnor4[305] = 1'b0 ^~ inbuffer_data[305];
assign xnor4[306] = 1'b1 ^~ inbuffer_data[306];
assign xnor4[307] = 1'b0 ^~ inbuffer_data[307];
assign xnor4[308] = 1'b1 ^~ inbuffer_data[308];
assign xnor4[309] = 1'b1 ^~ inbuffer_data[309];
assign xnor4[310] = 1'b0 ^~ inbuffer_data[310];
assign xnor4[311] = 1'b0 ^~ inbuffer_data[311];
assign xnor4[312] = 1'b0 ^~ inbuffer_data[312];
assign xnor4[313] = 1'b1 ^~ inbuffer_data[313];
assign xnor4[314] = 1'b1 ^~ inbuffer_data[314];
assign xnor4[315] = 1'b1 ^~ inbuffer_data[315];
assign xnor4[316] = 1'b1 ^~ inbuffer_data[316];
assign xnor4[317] = 1'b1 ^~ inbuffer_data[317];
assign xnor4[318] = 1'b1 ^~ inbuffer_data[318];
assign xnor4[319] = 1'b1 ^~ inbuffer_data[319];
assign xnor4[320] = 1'b1 ^~ inbuffer_data[320];
assign xnor4[321] = 1'b0 ^~ inbuffer_data[321];
assign xnor4[322] = 1'b0 ^~ inbuffer_data[322];
assign xnor4[323] = 1'b1 ^~ inbuffer_data[323];
assign xnor4[324] = 1'b1 ^~ inbuffer_data[324];
assign xnor4[325] = 1'b1 ^~ inbuffer_data[325];
assign xnor4[326] = 1'b0 ^~ inbuffer_data[326];
assign xnor4[327] = 1'b1 ^~ inbuffer_data[327];
assign xnor4[328] = 1'b0 ^~ inbuffer_data[328];
assign xnor4[329] = 1'b1 ^~ inbuffer_data[329];
assign xnor4[330] = 1'b0 ^~ inbuffer_data[330];
assign xnor4[331] = 1'b0 ^~ inbuffer_data[331];
assign xnor4[332] = 1'b0 ^~ inbuffer_data[332];
assign xnor4[333] = 1'b0 ^~ inbuffer_data[333];
assign xnor4[334] = 1'b0 ^~ inbuffer_data[334];
assign xnor4[335] = 1'b1 ^~ inbuffer_data[335];
assign xnor4[336] = 1'b1 ^~ inbuffer_data[336];
assign xnor4[337] = 1'b1 ^~ inbuffer_data[337];
assign xnor4[338] = 1'b0 ^~ inbuffer_data[338];
assign xnor4[339] = 1'b0 ^~ inbuffer_data[339];
assign xnor4[340] = 1'b0 ^~ inbuffer_data[340];
assign xnor4[341] = 1'b0 ^~ inbuffer_data[341];
assign xnor4[342] = 1'b1 ^~ inbuffer_data[342];
assign xnor4[343] = 1'b1 ^~ inbuffer_data[343];
assign xnor4[344] = 1'b1 ^~ inbuffer_data[344];
assign xnor4[345] = 1'b1 ^~ inbuffer_data[345];
assign xnor4[346] = 1'b1 ^~ inbuffer_data[346];
assign xnor4[347] = 1'b1 ^~ inbuffer_data[347];
assign xnor4[348] = 1'b1 ^~ inbuffer_data[348];
assign xnor4[349] = 1'b1 ^~ inbuffer_data[349];
assign xnor4[350] = 1'b0 ^~ inbuffer_data[350];
assign xnor4[351] = 1'b0 ^~ inbuffer_data[351];
assign xnor4[352] = 1'b1 ^~ inbuffer_data[352];
assign xnor4[353] = 1'b1 ^~ inbuffer_data[353];
assign xnor4[354] = 1'b1 ^~ inbuffer_data[354];
assign xnor4[355] = 1'b0 ^~ inbuffer_data[355];
assign xnor4[356] = 1'b0 ^~ inbuffer_data[356];
assign xnor4[357] = 1'b1 ^~ inbuffer_data[357];
assign xnor4[358] = 1'b1 ^~ inbuffer_data[358];
assign xnor4[359] = 1'b0 ^~ inbuffer_data[359];
assign xnor4[360] = 1'b0 ^~ inbuffer_data[360];
assign xnor4[361] = 1'b1 ^~ inbuffer_data[361];
assign xnor4[362] = 1'b0 ^~ inbuffer_data[362];
assign xnor4[363] = 1'b1 ^~ inbuffer_data[363];
assign xnor4[364] = 1'b0 ^~ inbuffer_data[364];
assign xnor4[365] = 1'b1 ^~ inbuffer_data[365];
assign xnor4[366] = 1'b0 ^~ inbuffer_data[366];
assign xnor4[367] = 1'b1 ^~ inbuffer_data[367];
assign xnor4[368] = 1'b0 ^~ inbuffer_data[368];
assign xnor4[369] = 1'b1 ^~ inbuffer_data[369];
assign xnor4[370] = 1'b1 ^~ inbuffer_data[370];
assign xnor4[371] = 1'b1 ^~ inbuffer_data[371];
assign xnor4[372] = 1'b1 ^~ inbuffer_data[372];
assign xnor4[373] = 1'b1 ^~ inbuffer_data[373];
assign xnor4[374] = 1'b1 ^~ inbuffer_data[374];
assign xnor4[375] = 1'b1 ^~ inbuffer_data[375];
assign xnor4[376] = 1'b1 ^~ inbuffer_data[376];
assign xnor4[377] = 1'b1 ^~ inbuffer_data[377];
assign xnor4[378] = 1'b0 ^~ inbuffer_data[378];
assign xnor4[379] = 1'b1 ^~ inbuffer_data[379];
assign xnor4[380] = 1'b1 ^~ inbuffer_data[380];
assign xnor4[381] = 1'b1 ^~ inbuffer_data[381];
assign xnor4[382] = 1'b1 ^~ inbuffer_data[382];
assign xnor4[383] = 1'b0 ^~ inbuffer_data[383];
assign xnor4[384] = 1'b1 ^~ inbuffer_data[384];
assign xnor4[385] = 1'b1 ^~ inbuffer_data[385];
assign xnor4[386] = 1'b1 ^~ inbuffer_data[386];
assign xnor4[387] = 1'b0 ^~ inbuffer_data[387];
assign xnor4[388] = 1'b0 ^~ inbuffer_data[388];
assign xnor4[389] = 1'b1 ^~ inbuffer_data[389];
assign xnor4[390] = 1'b0 ^~ inbuffer_data[390];
assign xnor4[391] = 1'b1 ^~ inbuffer_data[391];
assign xnor4[392] = 1'b1 ^~ inbuffer_data[392];
assign xnor4[393] = 1'b0 ^~ inbuffer_data[393];
assign xnor4[394] = 1'b0 ^~ inbuffer_data[394];
assign xnor4[395] = 1'b0 ^~ inbuffer_data[395];
assign xnor4[396] = 1'b1 ^~ inbuffer_data[396];
assign xnor4[397] = 1'b1 ^~ inbuffer_data[397];
assign xnor4[398] = 1'b1 ^~ inbuffer_data[398];
assign xnor4[399] = 1'b1 ^~ inbuffer_data[399];
assign xnor4[400] = 1'b1 ^~ inbuffer_data[400];
assign xnor4[401] = 1'b1 ^~ inbuffer_data[401];
assign xnor4[402] = 1'b1 ^~ inbuffer_data[402];
assign xnor4[403] = 1'b1 ^~ inbuffer_data[403];
assign xnor4[404] = 1'b1 ^~ inbuffer_data[404];
assign xnor4[405] = 1'b1 ^~ inbuffer_data[405];
assign xnor4[406] = 1'b0 ^~ inbuffer_data[406];
assign xnor4[407] = 1'b1 ^~ inbuffer_data[407];
assign xnor4[408] = 1'b1 ^~ inbuffer_data[408];
assign xnor4[409] = 1'b1 ^~ inbuffer_data[409];
assign xnor4[410] = 1'b1 ^~ inbuffer_data[410];
assign xnor4[411] = 1'b1 ^~ inbuffer_data[411];
assign xnor4[412] = 1'b1 ^~ inbuffer_data[412];
assign xnor4[413] = 1'b1 ^~ inbuffer_data[413];
assign xnor4[414] = 1'b1 ^~ inbuffer_data[414];
assign xnor4[415] = 1'b0 ^~ inbuffer_data[415];
assign xnor4[416] = 1'b0 ^~ inbuffer_data[416];
assign xnor4[417] = 1'b1 ^~ inbuffer_data[417];
assign xnor4[418] = 1'b1 ^~ inbuffer_data[418];
assign xnor4[419] = 1'b1 ^~ inbuffer_data[419];
assign xnor4[420] = 1'b0 ^~ inbuffer_data[420];
assign xnor4[421] = 1'b1 ^~ inbuffer_data[421];
assign xnor4[422] = 1'b1 ^~ inbuffer_data[422];
assign xnor4[423] = 1'b1 ^~ inbuffer_data[423];
assign xnor4[424] = 1'b1 ^~ inbuffer_data[424];
assign xnor4[425] = 1'b1 ^~ inbuffer_data[425];
assign xnor4[426] = 1'b1 ^~ inbuffer_data[426];
assign xnor4[427] = 1'b1 ^~ inbuffer_data[427];
assign xnor4[428] = 1'b1 ^~ inbuffer_data[428];
assign xnor4[429] = 1'b1 ^~ inbuffer_data[429];
assign xnor4[430] = 1'b1 ^~ inbuffer_data[430];
assign xnor4[431] = 1'b1 ^~ inbuffer_data[431];
assign xnor4[432] = 1'b1 ^~ inbuffer_data[432];
assign xnor4[433] = 1'b0 ^~ inbuffer_data[433];
assign xnor4[434] = 1'b1 ^~ inbuffer_data[434];
assign xnor4[435] = 1'b1 ^~ inbuffer_data[435];
assign xnor4[436] = 1'b1 ^~ inbuffer_data[436];
assign xnor4[437] = 1'b1 ^~ inbuffer_data[437];
assign xnor4[438] = 1'b1 ^~ inbuffer_data[438];
assign xnor4[439] = 1'b1 ^~ inbuffer_data[439];
assign xnor4[440] = 1'b1 ^~ inbuffer_data[440];
assign xnor4[441] = 1'b0 ^~ inbuffer_data[441];
assign xnor4[442] = 1'b1 ^~ inbuffer_data[442];
assign xnor4[443] = 1'b0 ^~ inbuffer_data[443];
assign xnor4[444] = 1'b0 ^~ inbuffer_data[444];
assign xnor4[445] = 1'b0 ^~ inbuffer_data[445];
assign xnor4[446] = 1'b1 ^~ inbuffer_data[446];
assign xnor4[447] = 1'b0 ^~ inbuffer_data[447];
assign xnor4[448] = 1'b0 ^~ inbuffer_data[448];
assign xnor4[449] = 1'b1 ^~ inbuffer_data[449];
assign xnor4[450] = 1'b0 ^~ inbuffer_data[450];
assign xnor4[451] = 1'b1 ^~ inbuffer_data[451];
assign xnor4[452] = 1'b0 ^~ inbuffer_data[452];
assign xnor4[453] = 1'b1 ^~ inbuffer_data[453];
assign xnor4[454] = 1'b1 ^~ inbuffer_data[454];
assign xnor4[455] = 1'b1 ^~ inbuffer_data[455];
assign xnor4[456] = 1'b1 ^~ inbuffer_data[456];
assign xnor4[457] = 1'b1 ^~ inbuffer_data[457];
assign xnor4[458] = 1'b1 ^~ inbuffer_data[458];
assign xnor4[459] = 1'b0 ^~ inbuffer_data[459];
assign xnor4[460] = 1'b1 ^~ inbuffer_data[460];
assign xnor4[461] = 1'b1 ^~ inbuffer_data[461];
assign xnor4[462] = 1'b1 ^~ inbuffer_data[462];
assign xnor4[463] = 1'b1 ^~ inbuffer_data[463];
assign xnor4[464] = 1'b1 ^~ inbuffer_data[464];
assign xnor4[465] = 1'b1 ^~ inbuffer_data[465];
assign xnor4[466] = 1'b1 ^~ inbuffer_data[466];
assign xnor4[467] = 1'b1 ^~ inbuffer_data[467];
assign xnor4[468] = 1'b1 ^~ inbuffer_data[468];
assign xnor4[469] = 1'b0 ^~ inbuffer_data[469];
assign xnor4[470] = 1'b0 ^~ inbuffer_data[470];
assign xnor4[471] = 1'b1 ^~ inbuffer_data[471];
assign xnor4[472] = 1'b0 ^~ inbuffer_data[472];
assign xnor4[473] = 1'b0 ^~ inbuffer_data[473];
assign xnor4[474] = 1'b0 ^~ inbuffer_data[474];
assign xnor4[475] = 1'b1 ^~ inbuffer_data[475];
assign xnor4[476] = 1'b1 ^~ inbuffer_data[476];
assign xnor4[477] = 1'b1 ^~ inbuffer_data[477];
assign xnor4[478] = 1'b1 ^~ inbuffer_data[478];
assign xnor4[479] = 1'b0 ^~ inbuffer_data[479];
assign xnor4[480] = 1'b0 ^~ inbuffer_data[480];
assign xnor4[481] = 1'b0 ^~ inbuffer_data[481];
assign xnor4[482] = 1'b0 ^~ inbuffer_data[482];
assign xnor4[483] = 1'b1 ^~ inbuffer_data[483];
assign xnor4[484] = 1'b1 ^~ inbuffer_data[484];
assign xnor4[485] = 1'b1 ^~ inbuffer_data[485];
assign xnor4[486] = 1'b0 ^~ inbuffer_data[486];
assign xnor4[487] = 1'b0 ^~ inbuffer_data[487];
assign xnor4[488] = 1'b1 ^~ inbuffer_data[488];
assign xnor4[489] = 1'b1 ^~ inbuffer_data[489];
assign xnor4[490] = 1'b1 ^~ inbuffer_data[490];
assign xnor4[491] = 1'b1 ^~ inbuffer_data[491];
assign xnor4[492] = 1'b1 ^~ inbuffer_data[492];
assign xnor4[493] = 1'b1 ^~ inbuffer_data[493];
assign xnor4[494] = 1'b1 ^~ inbuffer_data[494];
assign xnor4[495] = 1'b0 ^~ inbuffer_data[495];
assign xnor4[496] = 1'b0 ^~ inbuffer_data[496];
assign xnor4[497] = 1'b0 ^~ inbuffer_data[497];
assign xnor4[498] = 1'b0 ^~ inbuffer_data[498];
assign xnor4[499] = 1'b0 ^~ inbuffer_data[499];
assign xnor4[500] = 1'b0 ^~ inbuffer_data[500];
assign xnor4[501] = 1'b0 ^~ inbuffer_data[501];
assign xnor4[502] = 1'b0 ^~ inbuffer_data[502];
assign xnor4[503] = 1'b0 ^~ inbuffer_data[503];
assign xnor4[504] = 1'b1 ^~ inbuffer_data[504];
assign xnor4[505] = 1'b0 ^~ inbuffer_data[505];
assign xnor4[506] = 1'b1 ^~ inbuffer_data[506];
assign xnor4[507] = 1'b0 ^~ inbuffer_data[507];
assign xnor4[508] = 1'b0 ^~ inbuffer_data[508];
assign xnor4[509] = 1'b0 ^~ inbuffer_data[509];
assign xnor4[510] = 1'b0 ^~ inbuffer_data[510];
assign xnor4[511] = 1'b1 ^~ inbuffer_data[511];
assign xnor4[512] = 1'b1 ^~ inbuffer_data[512];
assign xnor4[513] = 1'b0 ^~ inbuffer_data[513];
assign xnor4[514] = 1'b0 ^~ inbuffer_data[514];
assign xnor4[515] = 1'b0 ^~ inbuffer_data[515];
assign xnor4[516] = 1'b1 ^~ inbuffer_data[516];
assign xnor4[517] = 1'b1 ^~ inbuffer_data[517];
assign xnor4[518] = 1'b1 ^~ inbuffer_data[518];
assign xnor4[519] = 1'b1 ^~ inbuffer_data[519];
assign xnor4[520] = 1'b1 ^~ inbuffer_data[520];
assign xnor4[521] = 1'b1 ^~ inbuffer_data[521];
assign xnor4[522] = 1'b0 ^~ inbuffer_data[522];
assign xnor4[523] = 1'b0 ^~ inbuffer_data[523];
assign xnor4[524] = 1'b1 ^~ inbuffer_data[524];
assign xnor4[525] = 1'b1 ^~ inbuffer_data[525];
assign xnor4[526] = 1'b0 ^~ inbuffer_data[526];
assign xnor4[527] = 1'b0 ^~ inbuffer_data[527];
assign xnor4[528] = 1'b0 ^~ inbuffer_data[528];
assign xnor4[529] = 1'b0 ^~ inbuffer_data[529];
assign xnor4[530] = 1'b0 ^~ inbuffer_data[530];
assign xnor4[531] = 1'b0 ^~ inbuffer_data[531];
assign xnor4[532] = 1'b0 ^~ inbuffer_data[532];
assign xnor4[533] = 1'b0 ^~ inbuffer_data[533];
assign xnor4[534] = 1'b0 ^~ inbuffer_data[534];
assign xnor4[535] = 1'b0 ^~ inbuffer_data[535];
assign xnor4[536] = 1'b0 ^~ inbuffer_data[536];
assign xnor4[537] = 1'b1 ^~ inbuffer_data[537];
assign xnor4[538] = 1'b0 ^~ inbuffer_data[538];
assign xnor4[539] = 1'b0 ^~ inbuffer_data[539];
assign xnor4[540] = 1'b0 ^~ inbuffer_data[540];
assign xnor4[541] = 1'b0 ^~ inbuffer_data[541];
assign xnor4[542] = 1'b0 ^~ inbuffer_data[542];
assign xnor4[543] = 1'b0 ^~ inbuffer_data[543];
assign xnor4[544] = 1'b0 ^~ inbuffer_data[544];
assign xnor4[545] = 1'b0 ^~ inbuffer_data[545];
assign xnor4[546] = 1'b1 ^~ inbuffer_data[546];
assign xnor4[547] = 1'b1 ^~ inbuffer_data[547];
assign xnor4[548] = 1'b0 ^~ inbuffer_data[548];
assign xnor4[549] = 1'b0 ^~ inbuffer_data[549];
assign xnor4[550] = 1'b0 ^~ inbuffer_data[550];
assign xnor4[551] = 1'b0 ^~ inbuffer_data[551];
assign xnor4[552] = 1'b0 ^~ inbuffer_data[552];
assign xnor4[553] = 1'b0 ^~ inbuffer_data[553];
assign xnor4[554] = 1'b0 ^~ inbuffer_data[554];
assign xnor4[555] = 1'b0 ^~ inbuffer_data[555];
assign xnor4[556] = 1'b0 ^~ inbuffer_data[556];
assign xnor4[557] = 1'b0 ^~ inbuffer_data[557];
assign xnor4[558] = 1'b1 ^~ inbuffer_data[558];
assign xnor4[559] = 1'b0 ^~ inbuffer_data[559];
assign xnor4[560] = 1'b1 ^~ inbuffer_data[560];
assign xnor4[561] = 1'b0 ^~ inbuffer_data[561];
assign xnor4[562] = 1'b0 ^~ inbuffer_data[562];
assign xnor4[563] = 1'b1 ^~ inbuffer_data[563];
assign xnor4[564] = 1'b1 ^~ inbuffer_data[564];
assign xnor4[565] = 1'b0 ^~ inbuffer_data[565];
assign xnor4[566] = 1'b0 ^~ inbuffer_data[566];
assign xnor4[567] = 1'b0 ^~ inbuffer_data[567];
assign xnor4[568] = 1'b0 ^~ inbuffer_data[568];
assign xnor4[569] = 1'b0 ^~ inbuffer_data[569];
assign xnor4[570] = 1'b0 ^~ inbuffer_data[570];
assign xnor4[571] = 1'b0 ^~ inbuffer_data[571];
assign xnor4[572] = 1'b0 ^~ inbuffer_data[572];
assign xnor4[573] = 1'b0 ^~ inbuffer_data[573];
assign xnor4[574] = 1'b0 ^~ inbuffer_data[574];
assign xnor4[575] = 1'b1 ^~ inbuffer_data[575];
assign xnor4[576] = 1'b1 ^~ inbuffer_data[576];
assign xnor4[577] = 1'b1 ^~ inbuffer_data[577];
assign xnor4[578] = 1'b0 ^~ inbuffer_data[578];
assign xnor4[579] = 1'b0 ^~ inbuffer_data[579];
assign xnor4[580] = 1'b1 ^~ inbuffer_data[580];
assign xnor4[581] = 1'b0 ^~ inbuffer_data[581];
assign xnor4[582] = 1'b0 ^~ inbuffer_data[582];
assign xnor4[583] = 1'b0 ^~ inbuffer_data[583];
assign xnor4[584] = 1'b0 ^~ inbuffer_data[584];
assign xnor4[585] = 1'b0 ^~ inbuffer_data[585];
assign xnor4[586] = 1'b0 ^~ inbuffer_data[586];
assign xnor4[587] = 1'b1 ^~ inbuffer_data[587];
assign xnor4[588] = 1'b0 ^~ inbuffer_data[588];
assign xnor4[589] = 1'b1 ^~ inbuffer_data[589];
assign xnor4[590] = 1'b1 ^~ inbuffer_data[590];
assign xnor4[591] = 1'b1 ^~ inbuffer_data[591];
assign xnor4[592] = 1'b0 ^~ inbuffer_data[592];
assign xnor4[593] = 1'b0 ^~ inbuffer_data[593];
assign xnor4[594] = 1'b0 ^~ inbuffer_data[594];
assign xnor4[595] = 1'b0 ^~ inbuffer_data[595];
assign xnor4[596] = 1'b0 ^~ inbuffer_data[596];
assign xnor4[597] = 1'b0 ^~ inbuffer_data[597];
assign xnor4[598] = 1'b0 ^~ inbuffer_data[598];
assign xnor4[599] = 1'b1 ^~ inbuffer_data[599];
assign xnor4[600] = 1'b0 ^~ inbuffer_data[600];
assign xnor4[601] = 1'b0 ^~ inbuffer_data[601];
assign xnor4[602] = 1'b0 ^~ inbuffer_data[602];
assign xnor4[603] = 1'b0 ^~ inbuffer_data[603];
assign xnor4[604] = 1'b0 ^~ inbuffer_data[604];
assign xnor4[605] = 1'b0 ^~ inbuffer_data[605];
assign xnor4[606] = 1'b1 ^~ inbuffer_data[606];
assign xnor4[607] = 1'b0 ^~ inbuffer_data[607];
assign xnor4[608] = 1'b1 ^~ inbuffer_data[608];
assign xnor4[609] = 1'b1 ^~ inbuffer_data[609];
assign xnor4[610] = 1'b1 ^~ inbuffer_data[610];
assign xnor4[611] = 1'b0 ^~ inbuffer_data[611];
assign xnor4[612] = 1'b0 ^~ inbuffer_data[612];
assign xnor4[613] = 1'b1 ^~ inbuffer_data[613];
assign xnor4[614] = 1'b0 ^~ inbuffer_data[614];
assign xnor4[615] = 1'b1 ^~ inbuffer_data[615];
assign xnor4[616] = 1'b1 ^~ inbuffer_data[616];
assign xnor4[617] = 1'b1 ^~ inbuffer_data[617];
assign xnor4[618] = 1'b0 ^~ inbuffer_data[618];
assign xnor4[619] = 1'b0 ^~ inbuffer_data[619];
assign xnor4[620] = 1'b0 ^~ inbuffer_data[620];
assign xnor4[621] = 1'b0 ^~ inbuffer_data[621];
assign xnor4[622] = 1'b0 ^~ inbuffer_data[622];
assign xnor4[623] = 1'b0 ^~ inbuffer_data[623];
assign xnor4[624] = 1'b0 ^~ inbuffer_data[624];
assign xnor4[625] = 1'b0 ^~ inbuffer_data[625];
assign xnor4[626] = 1'b0 ^~ inbuffer_data[626];
assign xnor4[627] = 1'b1 ^~ inbuffer_data[627];
assign xnor4[628] = 1'b0 ^~ inbuffer_data[628];
assign xnor4[629] = 1'b0 ^~ inbuffer_data[629];
assign xnor4[630] = 1'b0 ^~ inbuffer_data[630];
assign xnor4[631] = 1'b1 ^~ inbuffer_data[631];
assign xnor4[632] = 1'b0 ^~ inbuffer_data[632];
assign xnor4[633] = 1'b1 ^~ inbuffer_data[633];
assign xnor4[634] = 1'b0 ^~ inbuffer_data[634];
assign xnor4[635] = 1'b1 ^~ inbuffer_data[635];
assign xnor4[636] = 1'b1 ^~ inbuffer_data[636];
assign xnor4[637] = 1'b1 ^~ inbuffer_data[637];
assign xnor4[638] = 1'b0 ^~ inbuffer_data[638];
assign xnor4[639] = 1'b1 ^~ inbuffer_data[639];
assign xnor4[640] = 1'b1 ^~ inbuffer_data[640];
assign xnor4[641] = 1'b1 ^~ inbuffer_data[641];
assign xnor4[642] = 1'b1 ^~ inbuffer_data[642];
assign xnor4[643] = 1'b1 ^~ inbuffer_data[643];
assign xnor4[644] = 1'b1 ^~ inbuffer_data[644];
assign xnor4[645] = 1'b0 ^~ inbuffer_data[645];
assign xnor4[646] = 1'b0 ^~ inbuffer_data[646];
assign xnor4[647] = 1'b0 ^~ inbuffer_data[647];
assign xnor4[648] = 1'b1 ^~ inbuffer_data[648];
assign xnor4[649] = 1'b0 ^~ inbuffer_data[649];
assign xnor4[650] = 1'b0 ^~ inbuffer_data[650];
assign xnor4[651] = 1'b0 ^~ inbuffer_data[651];
assign xnor4[652] = 1'b0 ^~ inbuffer_data[652];
assign xnor4[653] = 1'b1 ^~ inbuffer_data[653];
assign xnor4[654] = 1'b0 ^~ inbuffer_data[654];
assign xnor4[655] = 1'b1 ^~ inbuffer_data[655];
assign xnor4[656] = 1'b0 ^~ inbuffer_data[656];
assign xnor4[657] = 1'b0 ^~ inbuffer_data[657];
assign xnor4[658] = 1'b0 ^~ inbuffer_data[658];
assign xnor4[659] = 1'b1 ^~ inbuffer_data[659];
assign xnor4[660] = 1'b1 ^~ inbuffer_data[660];
assign xnor4[661] = 1'b1 ^~ inbuffer_data[661];
assign xnor4[662] = 1'b1 ^~ inbuffer_data[662];
assign xnor4[663] = 1'b1 ^~ inbuffer_data[663];
assign xnor4[664] = 1'b1 ^~ inbuffer_data[664];
assign xnor4[665] = 1'b1 ^~ inbuffer_data[665];
assign xnor4[666] = 1'b1 ^~ inbuffer_data[666];
assign xnor4[667] = 1'b1 ^~ inbuffer_data[667];
assign xnor4[668] = 1'b0 ^~ inbuffer_data[668];
assign xnor4[669] = 1'b0 ^~ inbuffer_data[669];
assign xnor4[670] = 1'b1 ^~ inbuffer_data[670];
assign xnor4[671] = 1'b1 ^~ inbuffer_data[671];
assign xnor4[672] = 1'b1 ^~ inbuffer_data[672];
assign xnor4[673] = 1'b1 ^~ inbuffer_data[673];
assign xnor4[674] = 1'b1 ^~ inbuffer_data[674];
assign xnor4[675] = 1'b1 ^~ inbuffer_data[675];
assign xnor4[676] = 1'b0 ^~ inbuffer_data[676];
assign xnor4[677] = 1'b1 ^~ inbuffer_data[677];
assign xnor4[678] = 1'b1 ^~ inbuffer_data[678];
assign xnor4[679] = 1'b1 ^~ inbuffer_data[679];
assign xnor4[680] = 1'b0 ^~ inbuffer_data[680];
assign xnor4[681] = 1'b1 ^~ inbuffer_data[681];
assign xnor4[682] = 1'b1 ^~ inbuffer_data[682];
assign xnor4[683] = 1'b1 ^~ inbuffer_data[683];
assign xnor4[684] = 1'b0 ^~ inbuffer_data[684];
assign xnor4[685] = 1'b0 ^~ inbuffer_data[685];
assign xnor4[686] = 1'b0 ^~ inbuffer_data[686];
assign xnor4[687] = 1'b0 ^~ inbuffer_data[687];
assign xnor4[688] = 1'b0 ^~ inbuffer_data[688];
assign xnor4[689] = 1'b0 ^~ inbuffer_data[689];
assign xnor4[690] = 1'b1 ^~ inbuffer_data[690];
assign xnor4[691] = 1'b1 ^~ inbuffer_data[691];
assign xnor4[692] = 1'b0 ^~ inbuffer_data[692];
assign xnor4[693] = 1'b0 ^~ inbuffer_data[693];
assign xnor4[694] = 1'b0 ^~ inbuffer_data[694];
assign xnor4[695] = 1'b1 ^~ inbuffer_data[695];
assign xnor4[696] = 1'b0 ^~ inbuffer_data[696];
assign xnor4[697] = 1'b1 ^~ inbuffer_data[697];
assign xnor4[698] = 1'b1 ^~ inbuffer_data[698];
assign xnor4[699] = 1'b1 ^~ inbuffer_data[699];
assign xnor4[700] = 1'b0 ^~ inbuffer_data[700];
assign xnor4[701] = 1'b1 ^~ inbuffer_data[701];
assign xnor4[702] = 1'b0 ^~ inbuffer_data[702];
assign xnor4[703] = 1'b1 ^~ inbuffer_data[703];
assign xnor4[704] = 1'b1 ^~ inbuffer_data[704];
assign xnor4[705] = 1'b0 ^~ inbuffer_data[705];
assign xnor4[706] = 1'b1 ^~ inbuffer_data[706];
assign xnor4[707] = 1'b0 ^~ inbuffer_data[707];
assign xnor4[708] = 1'b0 ^~ inbuffer_data[708];
assign xnor4[709] = 1'b0 ^~ inbuffer_data[709];
assign xnor4[710] = 1'b0 ^~ inbuffer_data[710];
assign xnor4[711] = 1'b0 ^~ inbuffer_data[711];
assign xnor4[712] = 1'b0 ^~ inbuffer_data[712];
assign xnor4[713] = 1'b0 ^~ inbuffer_data[713];
assign xnor4[714] = 1'b0 ^~ inbuffer_data[714];
assign xnor4[715] = 1'b0 ^~ inbuffer_data[715];
assign xnor4[716] = 1'b0 ^~ inbuffer_data[716];
assign xnor4[717] = 1'b0 ^~ inbuffer_data[717];
assign xnor4[718] = 1'b0 ^~ inbuffer_data[718];
assign xnor4[719] = 1'b0 ^~ inbuffer_data[719];
assign xnor4[720] = 1'b0 ^~ inbuffer_data[720];
assign xnor4[721] = 1'b0 ^~ inbuffer_data[721];
assign xnor4[722] = 1'b1 ^~ inbuffer_data[722];
assign xnor4[723] = 1'b0 ^~ inbuffer_data[723];
assign xnor4[724] = 1'b1 ^~ inbuffer_data[724];
assign xnor4[725] = 1'b1 ^~ inbuffer_data[725];
assign xnor4[726] = 1'b0 ^~ inbuffer_data[726];
assign xnor4[727] = 1'b1 ^~ inbuffer_data[727];
assign xnor4[728] = 1'b1 ^~ inbuffer_data[728];
assign xnor4[729] = 1'b0 ^~ inbuffer_data[729];
assign xnor4[730] = 1'b0 ^~ inbuffer_data[730];
assign xnor4[731] = 1'b1 ^~ inbuffer_data[731];
assign xnor4[732] = 1'b1 ^~ inbuffer_data[732];
assign xnor4[733] = 1'b1 ^~ inbuffer_data[733];
assign xnor4[734] = 1'b0 ^~ inbuffer_data[734];
assign xnor4[735] = 1'b0 ^~ inbuffer_data[735];
assign xnor4[736] = 1'b0 ^~ inbuffer_data[736];
assign xnor4[737] = 1'b0 ^~ inbuffer_data[737];
assign xnor4[738] = 1'b0 ^~ inbuffer_data[738];
assign xnor4[739] = 1'b0 ^~ inbuffer_data[739];
assign xnor4[740] = 1'b0 ^~ inbuffer_data[740];
assign xnor4[741] = 1'b0 ^~ inbuffer_data[741];
assign xnor4[742] = 1'b0 ^~ inbuffer_data[742];
assign xnor4[743] = 1'b0 ^~ inbuffer_data[743];
assign xnor4[744] = 1'b0 ^~ inbuffer_data[744];
assign xnor4[745] = 1'b0 ^~ inbuffer_data[745];
assign xnor4[746] = 1'b0 ^~ inbuffer_data[746];
assign xnor4[747] = 1'b0 ^~ inbuffer_data[747];
assign xnor4[748] = 1'b0 ^~ inbuffer_data[748];
assign xnor4[749] = 1'b1 ^~ inbuffer_data[749];
assign xnor4[750] = 1'b0 ^~ inbuffer_data[750];
assign xnor4[751] = 1'b1 ^~ inbuffer_data[751];
assign xnor4[752] = 1'b1 ^~ inbuffer_data[752];
assign xnor4[753] = 1'b0 ^~ inbuffer_data[753];
assign xnor4[754] = 1'b1 ^~ inbuffer_data[754];
assign xnor4[755] = 1'b1 ^~ inbuffer_data[755];
assign xnor4[756] = 1'b0 ^~ inbuffer_data[756];
assign xnor4[757] = 1'b1 ^~ inbuffer_data[757];
assign xnor4[758] = 1'b0 ^~ inbuffer_data[758];
assign xnor4[759] = 1'b0 ^~ inbuffer_data[759];
assign xnor4[760] = 1'b0 ^~ inbuffer_data[760];
assign xnor4[761] = 1'b1 ^~ inbuffer_data[761];
assign xnor4[762] = 1'b1 ^~ inbuffer_data[762];
assign xnor4[763] = 1'b0 ^~ inbuffer_data[763];
assign xnor4[764] = 1'b0 ^~ inbuffer_data[764];
assign xnor4[765] = 1'b1 ^~ inbuffer_data[765];
assign xnor4[766] = 1'b0 ^~ inbuffer_data[766];
assign xnor4[767] = 1'b0 ^~ inbuffer_data[767];
assign xnor4[768] = 1'b0 ^~ inbuffer_data[768];
assign xnor4[769] = 1'b1 ^~ inbuffer_data[769];
assign xnor4[770] = 1'b1 ^~ inbuffer_data[770];
assign xnor4[771] = 1'b1 ^~ inbuffer_data[771];
assign xnor4[772] = 1'b1 ^~ inbuffer_data[772];
assign xnor4[773] = 1'b1 ^~ inbuffer_data[773];
assign xnor4[774] = 1'b0 ^~ inbuffer_data[774];
assign xnor4[775] = 1'b1 ^~ inbuffer_data[775];
assign xnor4[776] = 1'b1 ^~ inbuffer_data[776];
assign xnor4[777] = 1'b0 ^~ inbuffer_data[777];
assign xnor4[778] = 1'b0 ^~ inbuffer_data[778];
assign xnor4[779] = 1'b1 ^~ inbuffer_data[779];
assign xnor4[780] = 1'b0 ^~ inbuffer_data[780];
assign xnor4[781] = 1'b1 ^~ inbuffer_data[781];
assign xnor4[782] = 1'b0 ^~ inbuffer_data[782];
assign xnor4[783] = 1'b0 ^~ inbuffer_data[783];
assign xnor5[0] = 1'b1 ^~ inbuffer_data[0];
assign xnor5[1] = 1'b1 ^~ inbuffer_data[1];
assign xnor5[2] = 1'b0 ^~ inbuffer_data[2];
assign xnor5[3] = 1'b0 ^~ inbuffer_data[3];
assign xnor5[4] = 1'b1 ^~ inbuffer_data[4];
assign xnor5[5] = 1'b1 ^~ inbuffer_data[5];
assign xnor5[6] = 1'b0 ^~ inbuffer_data[6];
assign xnor5[7] = 1'b0 ^~ inbuffer_data[7];
assign xnor5[8] = 1'b1 ^~ inbuffer_data[8];
assign xnor5[9] = 1'b0 ^~ inbuffer_data[9];
assign xnor5[10] = 1'b1 ^~ inbuffer_data[10];
assign xnor5[11] = 1'b1 ^~ inbuffer_data[11];
assign xnor5[12] = 1'b0 ^~ inbuffer_data[12];
assign xnor5[13] = 1'b0 ^~ inbuffer_data[13];
assign xnor5[14] = 1'b1 ^~ inbuffer_data[14];
assign xnor5[15] = 1'b0 ^~ inbuffer_data[15];
assign xnor5[16] = 1'b0 ^~ inbuffer_data[16];
assign xnor5[17] = 1'b0 ^~ inbuffer_data[17];
assign xnor5[18] = 1'b0 ^~ inbuffer_data[18];
assign xnor5[19] = 1'b1 ^~ inbuffer_data[19];
assign xnor5[20] = 1'b0 ^~ inbuffer_data[20];
assign xnor5[21] = 1'b1 ^~ inbuffer_data[21];
assign xnor5[22] = 1'b0 ^~ inbuffer_data[22];
assign xnor5[23] = 1'b1 ^~ inbuffer_data[23];
assign xnor5[24] = 1'b0 ^~ inbuffer_data[24];
assign xnor5[25] = 1'b0 ^~ inbuffer_data[25];
assign xnor5[26] = 1'b0 ^~ inbuffer_data[26];
assign xnor5[27] = 1'b1 ^~ inbuffer_data[27];
assign xnor5[28] = 1'b0 ^~ inbuffer_data[28];
assign xnor5[29] = 1'b0 ^~ inbuffer_data[29];
assign xnor5[30] = 1'b1 ^~ inbuffer_data[30];
assign xnor5[31] = 1'b1 ^~ inbuffer_data[31];
assign xnor5[32] = 1'b1 ^~ inbuffer_data[32];
assign xnor5[33] = 1'b0 ^~ inbuffer_data[33];
assign xnor5[34] = 1'b1 ^~ inbuffer_data[34];
assign xnor5[35] = 1'b0 ^~ inbuffer_data[35];
assign xnor5[36] = 1'b0 ^~ inbuffer_data[36];
assign xnor5[37] = 1'b1 ^~ inbuffer_data[37];
assign xnor5[38] = 1'b1 ^~ inbuffer_data[38];
assign xnor5[39] = 1'b1 ^~ inbuffer_data[39];
assign xnor5[40] = 1'b1 ^~ inbuffer_data[40];
assign xnor5[41] = 1'b1 ^~ inbuffer_data[41];
assign xnor5[42] = 1'b1 ^~ inbuffer_data[42];
assign xnor5[43] = 1'b0 ^~ inbuffer_data[43];
assign xnor5[44] = 1'b1 ^~ inbuffer_data[44];
assign xnor5[45] = 1'b0 ^~ inbuffer_data[45];
assign xnor5[46] = 1'b0 ^~ inbuffer_data[46];
assign xnor5[47] = 1'b1 ^~ inbuffer_data[47];
assign xnor5[48] = 1'b0 ^~ inbuffer_data[48];
assign xnor5[49] = 1'b1 ^~ inbuffer_data[49];
assign xnor5[50] = 1'b1 ^~ inbuffer_data[50];
assign xnor5[51] = 1'b1 ^~ inbuffer_data[51];
assign xnor5[52] = 1'b1 ^~ inbuffer_data[52];
assign xnor5[53] = 1'b0 ^~ inbuffer_data[53];
assign xnor5[54] = 1'b1 ^~ inbuffer_data[54];
assign xnor5[55] = 1'b0 ^~ inbuffer_data[55];
assign xnor5[56] = 1'b0 ^~ inbuffer_data[56];
assign xnor5[57] = 1'b1 ^~ inbuffer_data[57];
assign xnor5[58] = 1'b0 ^~ inbuffer_data[58];
assign xnor5[59] = 1'b0 ^~ inbuffer_data[59];
assign xnor5[60] = 1'b1 ^~ inbuffer_data[60];
assign xnor5[61] = 1'b1 ^~ inbuffer_data[61];
assign xnor5[62] = 1'b0 ^~ inbuffer_data[62];
assign xnor5[63] = 1'b0 ^~ inbuffer_data[63];
assign xnor5[64] = 1'b0 ^~ inbuffer_data[64];
assign xnor5[65] = 1'b1 ^~ inbuffer_data[65];
assign xnor5[66] = 1'b0 ^~ inbuffer_data[66];
assign xnor5[67] = 1'b0 ^~ inbuffer_data[67];
assign xnor5[68] = 1'b0 ^~ inbuffer_data[68];
assign xnor5[69] = 1'b1 ^~ inbuffer_data[69];
assign xnor5[70] = 1'b0 ^~ inbuffer_data[70];
assign xnor5[71] = 1'b0 ^~ inbuffer_data[71];
assign xnor5[72] = 1'b0 ^~ inbuffer_data[72];
assign xnor5[73] = 1'b0 ^~ inbuffer_data[73];
assign xnor5[74] = 1'b1 ^~ inbuffer_data[74];
assign xnor5[75] = 1'b1 ^~ inbuffer_data[75];
assign xnor5[76] = 1'b0 ^~ inbuffer_data[76];
assign xnor5[77] = 1'b0 ^~ inbuffer_data[77];
assign xnor5[78] = 1'b0 ^~ inbuffer_data[78];
assign xnor5[79] = 1'b0 ^~ inbuffer_data[79];
assign xnor5[80] = 1'b0 ^~ inbuffer_data[80];
assign xnor5[81] = 1'b0 ^~ inbuffer_data[81];
assign xnor5[82] = 1'b0 ^~ inbuffer_data[82];
assign xnor5[83] = 1'b0 ^~ inbuffer_data[83];
assign xnor5[84] = 1'b1 ^~ inbuffer_data[84];
assign xnor5[85] = 1'b0 ^~ inbuffer_data[85];
assign xnor5[86] = 1'b0 ^~ inbuffer_data[86];
assign xnor5[87] = 1'b1 ^~ inbuffer_data[87];
assign xnor5[88] = 1'b1 ^~ inbuffer_data[88];
assign xnor5[89] = 1'b0 ^~ inbuffer_data[89];
assign xnor5[90] = 1'b1 ^~ inbuffer_data[90];
assign xnor5[91] = 1'b0 ^~ inbuffer_data[91];
assign xnor5[92] = 1'b0 ^~ inbuffer_data[92];
assign xnor5[93] = 1'b1 ^~ inbuffer_data[93];
assign xnor5[94] = 1'b0 ^~ inbuffer_data[94];
assign xnor5[95] = 1'b0 ^~ inbuffer_data[95];
assign xnor5[96] = 1'b0 ^~ inbuffer_data[96];
assign xnor5[97] = 1'b0 ^~ inbuffer_data[97];
assign xnor5[98] = 1'b0 ^~ inbuffer_data[98];
assign xnor5[99] = 1'b0 ^~ inbuffer_data[99];
assign xnor5[100] = 1'b0 ^~ inbuffer_data[100];
assign xnor5[101] = 1'b0 ^~ inbuffer_data[101];
assign xnor5[102] = 1'b0 ^~ inbuffer_data[102];
assign xnor5[103] = 1'b0 ^~ inbuffer_data[103];
assign xnor5[104] = 1'b1 ^~ inbuffer_data[104];
assign xnor5[105] = 1'b1 ^~ inbuffer_data[105];
assign xnor5[106] = 1'b1 ^~ inbuffer_data[106];
assign xnor5[107] = 1'b0 ^~ inbuffer_data[107];
assign xnor5[108] = 1'b0 ^~ inbuffer_data[108];
assign xnor5[109] = 1'b1 ^~ inbuffer_data[109];
assign xnor5[110] = 1'b0 ^~ inbuffer_data[110];
assign xnor5[111] = 1'b0 ^~ inbuffer_data[111];
assign xnor5[112] = 1'b1 ^~ inbuffer_data[112];
assign xnor5[113] = 1'b0 ^~ inbuffer_data[113];
assign xnor5[114] = 1'b0 ^~ inbuffer_data[114];
assign xnor5[115] = 1'b0 ^~ inbuffer_data[115];
assign xnor5[116] = 1'b1 ^~ inbuffer_data[116];
assign xnor5[117] = 1'b0 ^~ inbuffer_data[117];
assign xnor5[118] = 1'b0 ^~ inbuffer_data[118];
assign xnor5[119] = 1'b0 ^~ inbuffer_data[119];
assign xnor5[120] = 1'b0 ^~ inbuffer_data[120];
assign xnor5[121] = 1'b0 ^~ inbuffer_data[121];
assign xnor5[122] = 1'b0 ^~ inbuffer_data[122];
assign xnor5[123] = 1'b0 ^~ inbuffer_data[123];
assign xnor5[124] = 1'b0 ^~ inbuffer_data[124];
assign xnor5[125] = 1'b0 ^~ inbuffer_data[125];
assign xnor5[126] = 1'b0 ^~ inbuffer_data[126];
assign xnor5[127] = 1'b1 ^~ inbuffer_data[127];
assign xnor5[128] = 1'b1 ^~ inbuffer_data[128];
assign xnor5[129] = 1'b0 ^~ inbuffer_data[129];
assign xnor5[130] = 1'b1 ^~ inbuffer_data[130];
assign xnor5[131] = 1'b1 ^~ inbuffer_data[131];
assign xnor5[132] = 1'b0 ^~ inbuffer_data[132];
assign xnor5[133] = 1'b1 ^~ inbuffer_data[133];
assign xnor5[134] = 1'b1 ^~ inbuffer_data[134];
assign xnor5[135] = 1'b0 ^~ inbuffer_data[135];
assign xnor5[136] = 1'b1 ^~ inbuffer_data[136];
assign xnor5[137] = 1'b1 ^~ inbuffer_data[137];
assign xnor5[138] = 1'b0 ^~ inbuffer_data[138];
assign xnor5[139] = 1'b0 ^~ inbuffer_data[139];
assign xnor5[140] = 1'b0 ^~ inbuffer_data[140];
assign xnor5[141] = 1'b1 ^~ inbuffer_data[141];
assign xnor5[142] = 1'b0 ^~ inbuffer_data[142];
assign xnor5[143] = 1'b1 ^~ inbuffer_data[143];
assign xnor5[144] = 1'b0 ^~ inbuffer_data[144];
assign xnor5[145] = 1'b0 ^~ inbuffer_data[145];
assign xnor5[146] = 1'b0 ^~ inbuffer_data[146];
assign xnor5[147] = 1'b0 ^~ inbuffer_data[147];
assign xnor5[148] = 1'b0 ^~ inbuffer_data[148];
assign xnor5[149] = 1'b1 ^~ inbuffer_data[149];
assign xnor5[150] = 1'b1 ^~ inbuffer_data[150];
assign xnor5[151] = 1'b0 ^~ inbuffer_data[151];
assign xnor5[152] = 1'b0 ^~ inbuffer_data[152];
assign xnor5[153] = 1'b1 ^~ inbuffer_data[153];
assign xnor5[154] = 1'b0 ^~ inbuffer_data[154];
assign xnor5[155] = 1'b0 ^~ inbuffer_data[155];
assign xnor5[156] = 1'b1 ^~ inbuffer_data[156];
assign xnor5[157] = 1'b1 ^~ inbuffer_data[157];
assign xnor5[158] = 1'b1 ^~ inbuffer_data[158];
assign xnor5[159] = 1'b0 ^~ inbuffer_data[159];
assign xnor5[160] = 1'b1 ^~ inbuffer_data[160];
assign xnor5[161] = 1'b1 ^~ inbuffer_data[161];
assign xnor5[162] = 1'b1 ^~ inbuffer_data[162];
assign xnor5[163] = 1'b1 ^~ inbuffer_data[163];
assign xnor5[164] = 1'b1 ^~ inbuffer_data[164];
assign xnor5[165] = 1'b1 ^~ inbuffer_data[165];
assign xnor5[166] = 1'b0 ^~ inbuffer_data[166];
assign xnor5[167] = 1'b0 ^~ inbuffer_data[167];
assign xnor5[168] = 1'b1 ^~ inbuffer_data[168];
assign xnor5[169] = 1'b0 ^~ inbuffer_data[169];
assign xnor5[170] = 1'b1 ^~ inbuffer_data[170];
assign xnor5[171] = 1'b0 ^~ inbuffer_data[171];
assign xnor5[172] = 1'b0 ^~ inbuffer_data[172];
assign xnor5[173] = 1'b0 ^~ inbuffer_data[173];
assign xnor5[174] = 1'b0 ^~ inbuffer_data[174];
assign xnor5[175] = 1'b1 ^~ inbuffer_data[175];
assign xnor5[176] = 1'b0 ^~ inbuffer_data[176];
assign xnor5[177] = 1'b0 ^~ inbuffer_data[177];
assign xnor5[178] = 1'b0 ^~ inbuffer_data[178];
assign xnor5[179] = 1'b0 ^~ inbuffer_data[179];
assign xnor5[180] = 1'b1 ^~ inbuffer_data[180];
assign xnor5[181] = 1'b0 ^~ inbuffer_data[181];
assign xnor5[182] = 1'b1 ^~ inbuffer_data[182];
assign xnor5[183] = 1'b0 ^~ inbuffer_data[183];
assign xnor5[184] = 1'b1 ^~ inbuffer_data[184];
assign xnor5[185] = 1'b1 ^~ inbuffer_data[185];
assign xnor5[186] = 1'b0 ^~ inbuffer_data[186];
assign xnor5[187] = 1'b1 ^~ inbuffer_data[187];
assign xnor5[188] = 1'b1 ^~ inbuffer_data[188];
assign xnor5[189] = 1'b1 ^~ inbuffer_data[189];
assign xnor5[190] = 1'b1 ^~ inbuffer_data[190];
assign xnor5[191] = 1'b1 ^~ inbuffer_data[191];
assign xnor5[192] = 1'b1 ^~ inbuffer_data[192];
assign xnor5[193] = 1'b1 ^~ inbuffer_data[193];
assign xnor5[194] = 1'b1 ^~ inbuffer_data[194];
assign xnor5[195] = 1'b0 ^~ inbuffer_data[195];
assign xnor5[196] = 1'b1 ^~ inbuffer_data[196];
assign xnor5[197] = 1'b0 ^~ inbuffer_data[197];
assign xnor5[198] = 1'b0 ^~ inbuffer_data[198];
assign xnor5[199] = 1'b1 ^~ inbuffer_data[199];
assign xnor5[200] = 1'b0 ^~ inbuffer_data[200];
assign xnor5[201] = 1'b0 ^~ inbuffer_data[201];
assign xnor5[202] = 1'b0 ^~ inbuffer_data[202];
assign xnor5[203] = 1'b0 ^~ inbuffer_data[203];
assign xnor5[204] = 1'b1 ^~ inbuffer_data[204];
assign xnor5[205] = 1'b0 ^~ inbuffer_data[205];
assign xnor5[206] = 1'b0 ^~ inbuffer_data[206];
assign xnor5[207] = 1'b1 ^~ inbuffer_data[207];
assign xnor5[208] = 1'b1 ^~ inbuffer_data[208];
assign xnor5[209] = 1'b0 ^~ inbuffer_data[209];
assign xnor5[210] = 1'b0 ^~ inbuffer_data[210];
assign xnor5[211] = 1'b1 ^~ inbuffer_data[211];
assign xnor5[212] = 1'b0 ^~ inbuffer_data[212];
assign xnor5[213] = 1'b0 ^~ inbuffer_data[213];
assign xnor5[214] = 1'b1 ^~ inbuffer_data[214];
assign xnor5[215] = 1'b0 ^~ inbuffer_data[215];
assign xnor5[216] = 1'b1 ^~ inbuffer_data[216];
assign xnor5[217] = 1'b1 ^~ inbuffer_data[217];
assign xnor5[218] = 1'b1 ^~ inbuffer_data[218];
assign xnor5[219] = 1'b1 ^~ inbuffer_data[219];
assign xnor5[220] = 1'b1 ^~ inbuffer_data[220];
assign xnor5[221] = 1'b1 ^~ inbuffer_data[221];
assign xnor5[222] = 1'b1 ^~ inbuffer_data[222];
assign xnor5[223] = 1'b0 ^~ inbuffer_data[223];
assign xnor5[224] = 1'b0 ^~ inbuffer_data[224];
assign xnor5[225] = 1'b1 ^~ inbuffer_data[225];
assign xnor5[226] = 1'b1 ^~ inbuffer_data[226];
assign xnor5[227] = 1'b0 ^~ inbuffer_data[227];
assign xnor5[228] = 1'b0 ^~ inbuffer_data[228];
assign xnor5[229] = 1'b0 ^~ inbuffer_data[229];
assign xnor5[230] = 1'b0 ^~ inbuffer_data[230];
assign xnor5[231] = 1'b1 ^~ inbuffer_data[231];
assign xnor5[232] = 1'b0 ^~ inbuffer_data[232];
assign xnor5[233] = 1'b0 ^~ inbuffer_data[233];
assign xnor5[234] = 1'b1 ^~ inbuffer_data[234];
assign xnor5[235] = 1'b1 ^~ inbuffer_data[235];
assign xnor5[236] = 1'b1 ^~ inbuffer_data[236];
assign xnor5[237] = 1'b0 ^~ inbuffer_data[237];
assign xnor5[238] = 1'b0 ^~ inbuffer_data[238];
assign xnor5[239] = 1'b0 ^~ inbuffer_data[239];
assign xnor5[240] = 1'b0 ^~ inbuffer_data[240];
assign xnor5[241] = 1'b1 ^~ inbuffer_data[241];
assign xnor5[242] = 1'b1 ^~ inbuffer_data[242];
assign xnor5[243] = 1'b1 ^~ inbuffer_data[243];
assign xnor5[244] = 1'b1 ^~ inbuffer_data[244];
assign xnor5[245] = 1'b1 ^~ inbuffer_data[245];
assign xnor5[246] = 1'b1 ^~ inbuffer_data[246];
assign xnor5[247] = 1'b1 ^~ inbuffer_data[247];
assign xnor5[248] = 1'b1 ^~ inbuffer_data[248];
assign xnor5[249] = 1'b1 ^~ inbuffer_data[249];
assign xnor5[250] = 1'b1 ^~ inbuffer_data[250];
assign xnor5[251] = 1'b0 ^~ inbuffer_data[251];
assign xnor5[252] = 1'b0 ^~ inbuffer_data[252];
assign xnor5[253] = 1'b0 ^~ inbuffer_data[253];
assign xnor5[254] = 1'b1 ^~ inbuffer_data[254];
assign xnor5[255] = 1'b0 ^~ inbuffer_data[255];
assign xnor5[256] = 1'b0 ^~ inbuffer_data[256];
assign xnor5[257] = 1'b0 ^~ inbuffer_data[257];
assign xnor5[258] = 1'b0 ^~ inbuffer_data[258];
assign xnor5[259] = 1'b0 ^~ inbuffer_data[259];
assign xnor5[260] = 1'b1 ^~ inbuffer_data[260];
assign xnor5[261] = 1'b0 ^~ inbuffer_data[261];
assign xnor5[262] = 1'b1 ^~ inbuffer_data[262];
assign xnor5[263] = 1'b1 ^~ inbuffer_data[263];
assign xnor5[264] = 1'b1 ^~ inbuffer_data[264];
assign xnor5[265] = 1'b0 ^~ inbuffer_data[265];
assign xnor5[266] = 1'b0 ^~ inbuffer_data[266];
assign xnor5[267] = 1'b0 ^~ inbuffer_data[267];
assign xnor5[268] = 1'b0 ^~ inbuffer_data[268];
assign xnor5[269] = 1'b0 ^~ inbuffer_data[269];
assign xnor5[270] = 1'b1 ^~ inbuffer_data[270];
assign xnor5[271] = 1'b0 ^~ inbuffer_data[271];
assign xnor5[272] = 1'b1 ^~ inbuffer_data[272];
assign xnor5[273] = 1'b1 ^~ inbuffer_data[273];
assign xnor5[274] = 1'b1 ^~ inbuffer_data[274];
assign xnor5[275] = 1'b1 ^~ inbuffer_data[275];
assign xnor5[276] = 1'b1 ^~ inbuffer_data[276];
assign xnor5[277] = 1'b1 ^~ inbuffer_data[277];
assign xnor5[278] = 1'b1 ^~ inbuffer_data[278];
assign xnor5[279] = 1'b0 ^~ inbuffer_data[279];
assign xnor5[280] = 1'b0 ^~ inbuffer_data[280];
assign xnor5[281] = 1'b1 ^~ inbuffer_data[281];
assign xnor5[282] = 1'b1 ^~ inbuffer_data[282];
assign xnor5[283] = 1'b1 ^~ inbuffer_data[283];
assign xnor5[284] = 1'b0 ^~ inbuffer_data[284];
assign xnor5[285] = 1'b0 ^~ inbuffer_data[285];
assign xnor5[286] = 1'b0 ^~ inbuffer_data[286];
assign xnor5[287] = 1'b1 ^~ inbuffer_data[287];
assign xnor5[288] = 1'b1 ^~ inbuffer_data[288];
assign xnor5[289] = 1'b1 ^~ inbuffer_data[289];
assign xnor5[290] = 1'b1 ^~ inbuffer_data[290];
assign xnor5[291] = 1'b1 ^~ inbuffer_data[291];
assign xnor5[292] = 1'b1 ^~ inbuffer_data[292];
assign xnor5[293] = 1'b1 ^~ inbuffer_data[293];
assign xnor5[294] = 1'b0 ^~ inbuffer_data[294];
assign xnor5[295] = 1'b0 ^~ inbuffer_data[295];
assign xnor5[296] = 1'b0 ^~ inbuffer_data[296];
assign xnor5[297] = 1'b0 ^~ inbuffer_data[297];
assign xnor5[298] = 1'b0 ^~ inbuffer_data[298];
assign xnor5[299] = 1'b0 ^~ inbuffer_data[299];
assign xnor5[300] = 1'b0 ^~ inbuffer_data[300];
assign xnor5[301] = 1'b1 ^~ inbuffer_data[301];
assign xnor5[302] = 1'b0 ^~ inbuffer_data[302];
assign xnor5[303] = 1'b1 ^~ inbuffer_data[303];
assign xnor5[304] = 1'b1 ^~ inbuffer_data[304];
assign xnor5[305] = 1'b1 ^~ inbuffer_data[305];
assign xnor5[306] = 1'b1 ^~ inbuffer_data[306];
assign xnor5[307] = 1'b1 ^~ inbuffer_data[307];
assign xnor5[308] = 1'b1 ^~ inbuffer_data[308];
assign xnor5[309] = 1'b0 ^~ inbuffer_data[309];
assign xnor5[310] = 1'b0 ^~ inbuffer_data[310];
assign xnor5[311] = 1'b0 ^~ inbuffer_data[311];
assign xnor5[312] = 1'b0 ^~ inbuffer_data[312];
assign xnor5[313] = 1'b0 ^~ inbuffer_data[313];
assign xnor5[314] = 1'b1 ^~ inbuffer_data[314];
assign xnor5[315] = 1'b1 ^~ inbuffer_data[315];
assign xnor5[316] = 1'b1 ^~ inbuffer_data[316];
assign xnor5[317] = 1'b1 ^~ inbuffer_data[317];
assign xnor5[318] = 1'b1 ^~ inbuffer_data[318];
assign xnor5[319] = 1'b1 ^~ inbuffer_data[319];
assign xnor5[320] = 1'b1 ^~ inbuffer_data[320];
assign xnor5[321] = 1'b1 ^~ inbuffer_data[321];
assign xnor5[322] = 1'b1 ^~ inbuffer_data[322];
assign xnor5[323] = 1'b0 ^~ inbuffer_data[323];
assign xnor5[324] = 1'b0 ^~ inbuffer_data[324];
assign xnor5[325] = 1'b0 ^~ inbuffer_data[325];
assign xnor5[326] = 1'b0 ^~ inbuffer_data[326];
assign xnor5[327] = 1'b0 ^~ inbuffer_data[327];
assign xnor5[328] = 1'b0 ^~ inbuffer_data[328];
assign xnor5[329] = 1'b0 ^~ inbuffer_data[329];
assign xnor5[330] = 1'b0 ^~ inbuffer_data[330];
assign xnor5[331] = 1'b0 ^~ inbuffer_data[331];
assign xnor5[332] = 1'b1 ^~ inbuffer_data[332];
assign xnor5[333] = 1'b1 ^~ inbuffer_data[333];
assign xnor5[334] = 1'b0 ^~ inbuffer_data[334];
assign xnor5[335] = 1'b1 ^~ inbuffer_data[335];
assign xnor5[336] = 1'b0 ^~ inbuffer_data[336];
assign xnor5[337] = 1'b0 ^~ inbuffer_data[337];
assign xnor5[338] = 1'b1 ^~ inbuffer_data[338];
assign xnor5[339] = 1'b0 ^~ inbuffer_data[339];
assign xnor5[340] = 1'b1 ^~ inbuffer_data[340];
assign xnor5[341] = 1'b1 ^~ inbuffer_data[341];
assign xnor5[342] = 1'b1 ^~ inbuffer_data[342];
assign xnor5[343] = 1'b1 ^~ inbuffer_data[343];
assign xnor5[344] = 1'b1 ^~ inbuffer_data[344];
assign xnor5[345] = 1'b1 ^~ inbuffer_data[345];
assign xnor5[346] = 1'b1 ^~ inbuffer_data[346];
assign xnor5[347] = 1'b1 ^~ inbuffer_data[347];
assign xnor5[348] = 1'b1 ^~ inbuffer_data[348];
assign xnor5[349] = 1'b1 ^~ inbuffer_data[349];
assign xnor5[350] = 1'b0 ^~ inbuffer_data[350];
assign xnor5[351] = 1'b1 ^~ inbuffer_data[351];
assign xnor5[352] = 1'b0 ^~ inbuffer_data[352];
assign xnor5[353] = 1'b0 ^~ inbuffer_data[353];
assign xnor5[354] = 1'b0 ^~ inbuffer_data[354];
assign xnor5[355] = 1'b0 ^~ inbuffer_data[355];
assign xnor5[356] = 1'b0 ^~ inbuffer_data[356];
assign xnor5[357] = 1'b0 ^~ inbuffer_data[357];
assign xnor5[358] = 1'b0 ^~ inbuffer_data[358];
assign xnor5[359] = 1'b0 ^~ inbuffer_data[359];
assign xnor5[360] = 1'b0 ^~ inbuffer_data[360];
assign xnor5[361] = 1'b1 ^~ inbuffer_data[361];
assign xnor5[362] = 1'b1 ^~ inbuffer_data[362];
assign xnor5[363] = 1'b0 ^~ inbuffer_data[363];
assign xnor5[364] = 1'b0 ^~ inbuffer_data[364];
assign xnor5[365] = 1'b1 ^~ inbuffer_data[365];
assign xnor5[366] = 1'b0 ^~ inbuffer_data[366];
assign xnor5[367] = 1'b0 ^~ inbuffer_data[367];
assign xnor5[368] = 1'b0 ^~ inbuffer_data[368];
assign xnor5[369] = 1'b1 ^~ inbuffer_data[369];
assign xnor5[370] = 1'b1 ^~ inbuffer_data[370];
assign xnor5[371] = 1'b1 ^~ inbuffer_data[371];
assign xnor5[372] = 1'b1 ^~ inbuffer_data[372];
assign xnor5[373] = 1'b0 ^~ inbuffer_data[373];
assign xnor5[374] = 1'b0 ^~ inbuffer_data[374];
assign xnor5[375] = 1'b1 ^~ inbuffer_data[375];
assign xnor5[376] = 1'b1 ^~ inbuffer_data[376];
assign xnor5[377] = 1'b1 ^~ inbuffer_data[377];
assign xnor5[378] = 1'b0 ^~ inbuffer_data[378];
assign xnor5[379] = 1'b0 ^~ inbuffer_data[379];
assign xnor5[380] = 1'b0 ^~ inbuffer_data[380];
assign xnor5[381] = 1'b0 ^~ inbuffer_data[381];
assign xnor5[382] = 1'b0 ^~ inbuffer_data[382];
assign xnor5[383] = 1'b1 ^~ inbuffer_data[383];
assign xnor5[384] = 1'b0 ^~ inbuffer_data[384];
assign xnor5[385] = 1'b0 ^~ inbuffer_data[385];
assign xnor5[386] = 1'b0 ^~ inbuffer_data[386];
assign xnor5[387] = 1'b0 ^~ inbuffer_data[387];
assign xnor5[388] = 1'b0 ^~ inbuffer_data[388];
assign xnor5[389] = 1'b0 ^~ inbuffer_data[389];
assign xnor5[390] = 1'b0 ^~ inbuffer_data[390];
assign xnor5[391] = 1'b0 ^~ inbuffer_data[391];
assign xnor5[392] = 1'b0 ^~ inbuffer_data[392];
assign xnor5[393] = 1'b1 ^~ inbuffer_data[393];
assign xnor5[394] = 1'b0 ^~ inbuffer_data[394];
assign xnor5[395] = 1'b0 ^~ inbuffer_data[395];
assign xnor5[396] = 1'b1 ^~ inbuffer_data[396];
assign xnor5[397] = 1'b0 ^~ inbuffer_data[397];
assign xnor5[398] = 1'b0 ^~ inbuffer_data[398];
assign xnor5[399] = 1'b0 ^~ inbuffer_data[399];
assign xnor5[400] = 1'b1 ^~ inbuffer_data[400];
assign xnor5[401] = 1'b1 ^~ inbuffer_data[401];
assign xnor5[402] = 1'b1 ^~ inbuffer_data[402];
assign xnor5[403] = 1'b1 ^~ inbuffer_data[403];
assign xnor5[404] = 1'b0 ^~ inbuffer_data[404];
assign xnor5[405] = 1'b1 ^~ inbuffer_data[405];
assign xnor5[406] = 1'b0 ^~ inbuffer_data[406];
assign xnor5[407] = 1'b0 ^~ inbuffer_data[407];
assign xnor5[408] = 1'b0 ^~ inbuffer_data[408];
assign xnor5[409] = 1'b0 ^~ inbuffer_data[409];
assign xnor5[410] = 1'b0 ^~ inbuffer_data[410];
assign xnor5[411] = 1'b0 ^~ inbuffer_data[411];
assign xnor5[412] = 1'b1 ^~ inbuffer_data[412];
assign xnor5[413] = 1'b0 ^~ inbuffer_data[413];
assign xnor5[414] = 1'b0 ^~ inbuffer_data[414];
assign xnor5[415] = 1'b0 ^~ inbuffer_data[415];
assign xnor5[416] = 1'b0 ^~ inbuffer_data[416];
assign xnor5[417] = 1'b1 ^~ inbuffer_data[417];
assign xnor5[418] = 1'b1 ^~ inbuffer_data[418];
assign xnor5[419] = 1'b0 ^~ inbuffer_data[419];
assign xnor5[420] = 1'b1 ^~ inbuffer_data[420];
assign xnor5[421] = 1'b1 ^~ inbuffer_data[421];
assign xnor5[422] = 1'b0 ^~ inbuffer_data[422];
assign xnor5[423] = 1'b0 ^~ inbuffer_data[423];
assign xnor5[424] = 1'b1 ^~ inbuffer_data[424];
assign xnor5[425] = 1'b0 ^~ inbuffer_data[425];
assign xnor5[426] = 1'b0 ^~ inbuffer_data[426];
assign xnor5[427] = 1'b0 ^~ inbuffer_data[427];
assign xnor5[428] = 1'b1 ^~ inbuffer_data[428];
assign xnor5[429] = 1'b1 ^~ inbuffer_data[429];
assign xnor5[430] = 1'b1 ^~ inbuffer_data[430];
assign xnor5[431] = 1'b1 ^~ inbuffer_data[431];
assign xnor5[432] = 1'b0 ^~ inbuffer_data[432];
assign xnor5[433] = 1'b1 ^~ inbuffer_data[433];
assign xnor5[434] = 1'b0 ^~ inbuffer_data[434];
assign xnor5[435] = 1'b0 ^~ inbuffer_data[435];
assign xnor5[436] = 1'b0 ^~ inbuffer_data[436];
assign xnor5[437] = 1'b0 ^~ inbuffer_data[437];
assign xnor5[438] = 1'b0 ^~ inbuffer_data[438];
assign xnor5[439] = 1'b0 ^~ inbuffer_data[439];
assign xnor5[440] = 1'b0 ^~ inbuffer_data[440];
assign xnor5[441] = 1'b0 ^~ inbuffer_data[441];
assign xnor5[442] = 1'b0 ^~ inbuffer_data[442];
assign xnor5[443] = 1'b0 ^~ inbuffer_data[443];
assign xnor5[444] = 1'b0 ^~ inbuffer_data[444];
assign xnor5[445] = 1'b0 ^~ inbuffer_data[445];
assign xnor5[446] = 1'b0 ^~ inbuffer_data[446];
assign xnor5[447] = 1'b0 ^~ inbuffer_data[447];
assign xnor5[448] = 1'b0 ^~ inbuffer_data[448];
assign xnor5[449] = 1'b0 ^~ inbuffer_data[449];
assign xnor5[450] = 1'b1 ^~ inbuffer_data[450];
assign xnor5[451] = 1'b0 ^~ inbuffer_data[451];
assign xnor5[452] = 1'b0 ^~ inbuffer_data[452];
assign xnor5[453] = 1'b0 ^~ inbuffer_data[453];
assign xnor5[454] = 1'b0 ^~ inbuffer_data[454];
assign xnor5[455] = 1'b0 ^~ inbuffer_data[455];
assign xnor5[456] = 1'b0 ^~ inbuffer_data[456];
assign xnor5[457] = 1'b0 ^~ inbuffer_data[457];
assign xnor5[458] = 1'b0 ^~ inbuffer_data[458];
assign xnor5[459] = 1'b0 ^~ inbuffer_data[459];
assign xnor5[460] = 1'b0 ^~ inbuffer_data[460];
assign xnor5[461] = 1'b0 ^~ inbuffer_data[461];
assign xnor5[462] = 1'b0 ^~ inbuffer_data[462];
assign xnor5[463] = 1'b0 ^~ inbuffer_data[463];
assign xnor5[464] = 1'b0 ^~ inbuffer_data[464];
assign xnor5[465] = 1'b0 ^~ inbuffer_data[465];
assign xnor5[466] = 1'b0 ^~ inbuffer_data[466];
assign xnor5[467] = 1'b0 ^~ inbuffer_data[467];
assign xnor5[468] = 1'b1 ^~ inbuffer_data[468];
assign xnor5[469] = 1'b0 ^~ inbuffer_data[469];
assign xnor5[470] = 1'b1 ^~ inbuffer_data[470];
assign xnor5[471] = 1'b0 ^~ inbuffer_data[471];
assign xnor5[472] = 1'b1 ^~ inbuffer_data[472];
assign xnor5[473] = 1'b0 ^~ inbuffer_data[473];
assign xnor5[474] = 1'b0 ^~ inbuffer_data[474];
assign xnor5[475] = 1'b0 ^~ inbuffer_data[475];
assign xnor5[476] = 1'b0 ^~ inbuffer_data[476];
assign xnor5[477] = 1'b1 ^~ inbuffer_data[477];
assign xnor5[478] = 1'b1 ^~ inbuffer_data[478];
assign xnor5[479] = 1'b0 ^~ inbuffer_data[479];
assign xnor5[480] = 1'b0 ^~ inbuffer_data[480];
assign xnor5[481] = 1'b1 ^~ inbuffer_data[481];
assign xnor5[482] = 1'b1 ^~ inbuffer_data[482];
assign xnor5[483] = 1'b0 ^~ inbuffer_data[483];
assign xnor5[484] = 1'b0 ^~ inbuffer_data[484];
assign xnor5[485] = 1'b0 ^~ inbuffer_data[485];
assign xnor5[486] = 1'b0 ^~ inbuffer_data[486];
assign xnor5[487] = 1'b0 ^~ inbuffer_data[487];
assign xnor5[488] = 1'b0 ^~ inbuffer_data[488];
assign xnor5[489] = 1'b0 ^~ inbuffer_data[489];
assign xnor5[490] = 1'b0 ^~ inbuffer_data[490];
assign xnor5[491] = 1'b1 ^~ inbuffer_data[491];
assign xnor5[492] = 1'b0 ^~ inbuffer_data[492];
assign xnor5[493] = 1'b1 ^~ inbuffer_data[493];
assign xnor5[494] = 1'b1 ^~ inbuffer_data[494];
assign xnor5[495] = 1'b0 ^~ inbuffer_data[495];
assign xnor5[496] = 1'b1 ^~ inbuffer_data[496];
assign xnor5[497] = 1'b0 ^~ inbuffer_data[497];
assign xnor5[498] = 1'b0 ^~ inbuffer_data[498];
assign xnor5[499] = 1'b1 ^~ inbuffer_data[499];
assign xnor5[500] = 1'b1 ^~ inbuffer_data[500];
assign xnor5[501] = 1'b0 ^~ inbuffer_data[501];
assign xnor5[502] = 1'b1 ^~ inbuffer_data[502];
assign xnor5[503] = 1'b0 ^~ inbuffer_data[503];
assign xnor5[504] = 1'b0 ^~ inbuffer_data[504];
assign xnor5[505] = 1'b0 ^~ inbuffer_data[505];
assign xnor5[506] = 1'b0 ^~ inbuffer_data[506];
assign xnor5[507] = 1'b1 ^~ inbuffer_data[507];
assign xnor5[508] = 1'b1 ^~ inbuffer_data[508];
assign xnor5[509] = 1'b1 ^~ inbuffer_data[509];
assign xnor5[510] = 1'b1 ^~ inbuffer_data[510];
assign xnor5[511] = 1'b1 ^~ inbuffer_data[511];
assign xnor5[512] = 1'b1 ^~ inbuffer_data[512];
assign xnor5[513] = 1'b0 ^~ inbuffer_data[513];
assign xnor5[514] = 1'b0 ^~ inbuffer_data[514];
assign xnor5[515] = 1'b0 ^~ inbuffer_data[515];
assign xnor5[516] = 1'b0 ^~ inbuffer_data[516];
assign xnor5[517] = 1'b0 ^~ inbuffer_data[517];
assign xnor5[518] = 1'b1 ^~ inbuffer_data[518];
assign xnor5[519] = 1'b0 ^~ inbuffer_data[519];
assign xnor5[520] = 1'b0 ^~ inbuffer_data[520];
assign xnor5[521] = 1'b0 ^~ inbuffer_data[521];
assign xnor5[522] = 1'b0 ^~ inbuffer_data[522];
assign xnor5[523] = 1'b1 ^~ inbuffer_data[523];
assign xnor5[524] = 1'b0 ^~ inbuffer_data[524];
assign xnor5[525] = 1'b1 ^~ inbuffer_data[525];
assign xnor5[526] = 1'b1 ^~ inbuffer_data[526];
assign xnor5[527] = 1'b1 ^~ inbuffer_data[527];
assign xnor5[528] = 1'b0 ^~ inbuffer_data[528];
assign xnor5[529] = 1'b0 ^~ inbuffer_data[529];
assign xnor5[530] = 1'b1 ^~ inbuffer_data[530];
assign xnor5[531] = 1'b0 ^~ inbuffer_data[531];
assign xnor5[532] = 1'b0 ^~ inbuffer_data[532];
assign xnor5[533] = 1'b0 ^~ inbuffer_data[533];
assign xnor5[534] = 1'b1 ^~ inbuffer_data[534];
assign xnor5[535] = 1'b1 ^~ inbuffer_data[535];
assign xnor5[536] = 1'b1 ^~ inbuffer_data[536];
assign xnor5[537] = 1'b1 ^~ inbuffer_data[537];
assign xnor5[538] = 1'b1 ^~ inbuffer_data[538];
assign xnor5[539] = 1'b1 ^~ inbuffer_data[539];
assign xnor5[540] = 1'b1 ^~ inbuffer_data[540];
assign xnor5[541] = 1'b1 ^~ inbuffer_data[541];
assign xnor5[542] = 1'b1 ^~ inbuffer_data[542];
assign xnor5[543] = 1'b0 ^~ inbuffer_data[543];
assign xnor5[544] = 1'b0 ^~ inbuffer_data[544];
assign xnor5[545] = 1'b1 ^~ inbuffer_data[545];
assign xnor5[546] = 1'b0 ^~ inbuffer_data[546];
assign xnor5[547] = 1'b1 ^~ inbuffer_data[547];
assign xnor5[548] = 1'b0 ^~ inbuffer_data[548];
assign xnor5[549] = 1'b0 ^~ inbuffer_data[549];
assign xnor5[550] = 1'b1 ^~ inbuffer_data[550];
assign xnor5[551] = 1'b1 ^~ inbuffer_data[551];
assign xnor5[552] = 1'b1 ^~ inbuffer_data[552];
assign xnor5[553] = 1'b1 ^~ inbuffer_data[553];
assign xnor5[554] = 1'b1 ^~ inbuffer_data[554];
assign xnor5[555] = 1'b1 ^~ inbuffer_data[555];
assign xnor5[556] = 1'b1 ^~ inbuffer_data[556];
assign xnor5[557] = 1'b1 ^~ inbuffer_data[557];
assign xnor5[558] = 1'b0 ^~ inbuffer_data[558];
assign xnor5[559] = 1'b1 ^~ inbuffer_data[559];
assign xnor5[560] = 1'b0 ^~ inbuffer_data[560];
assign xnor5[561] = 1'b1 ^~ inbuffer_data[561];
assign xnor5[562] = 1'b0 ^~ inbuffer_data[562];
assign xnor5[563] = 1'b0 ^~ inbuffer_data[563];
assign xnor5[564] = 1'b0 ^~ inbuffer_data[564];
assign xnor5[565] = 1'b1 ^~ inbuffer_data[565];
assign xnor5[566] = 1'b1 ^~ inbuffer_data[566];
assign xnor5[567] = 1'b1 ^~ inbuffer_data[567];
assign xnor5[568] = 1'b1 ^~ inbuffer_data[568];
assign xnor5[569] = 1'b1 ^~ inbuffer_data[569];
assign xnor5[570] = 1'b1 ^~ inbuffer_data[570];
assign xnor5[571] = 1'b1 ^~ inbuffer_data[571];
assign xnor5[572] = 1'b1 ^~ inbuffer_data[572];
assign xnor5[573] = 1'b0 ^~ inbuffer_data[573];
assign xnor5[574] = 1'b0 ^~ inbuffer_data[574];
assign xnor5[575] = 1'b0 ^~ inbuffer_data[575];
assign xnor5[576] = 1'b1 ^~ inbuffer_data[576];
assign xnor5[577] = 1'b1 ^~ inbuffer_data[577];
assign xnor5[578] = 1'b1 ^~ inbuffer_data[578];
assign xnor5[579] = 1'b1 ^~ inbuffer_data[579];
assign xnor5[580] = 1'b1 ^~ inbuffer_data[580];
assign xnor5[581] = 1'b1 ^~ inbuffer_data[581];
assign xnor5[582] = 1'b1 ^~ inbuffer_data[582];
assign xnor5[583] = 1'b1 ^~ inbuffer_data[583];
assign xnor5[584] = 1'b0 ^~ inbuffer_data[584];
assign xnor5[585] = 1'b1 ^~ inbuffer_data[585];
assign xnor5[586] = 1'b0 ^~ inbuffer_data[586];
assign xnor5[587] = 1'b0 ^~ inbuffer_data[587];
assign xnor5[588] = 1'b0 ^~ inbuffer_data[588];
assign xnor5[589] = 1'b1 ^~ inbuffer_data[589];
assign xnor5[590] = 1'b1 ^~ inbuffer_data[590];
assign xnor5[591] = 1'b1 ^~ inbuffer_data[591];
assign xnor5[592] = 1'b0 ^~ inbuffer_data[592];
assign xnor5[593] = 1'b0 ^~ inbuffer_data[593];
assign xnor5[594] = 1'b1 ^~ inbuffer_data[594];
assign xnor5[595] = 1'b1 ^~ inbuffer_data[595];
assign xnor5[596] = 1'b1 ^~ inbuffer_data[596];
assign xnor5[597] = 1'b1 ^~ inbuffer_data[597];
assign xnor5[598] = 1'b1 ^~ inbuffer_data[598];
assign xnor5[599] = 1'b0 ^~ inbuffer_data[599];
assign xnor5[600] = 1'b1 ^~ inbuffer_data[600];
assign xnor5[601] = 1'b0 ^~ inbuffer_data[601];
assign xnor5[602] = 1'b1 ^~ inbuffer_data[602];
assign xnor5[603] = 1'b0 ^~ inbuffer_data[603];
assign xnor5[604] = 1'b0 ^~ inbuffer_data[604];
assign xnor5[605] = 1'b0 ^~ inbuffer_data[605];
assign xnor5[606] = 1'b1 ^~ inbuffer_data[606];
assign xnor5[607] = 1'b1 ^~ inbuffer_data[607];
assign xnor5[608] = 1'b1 ^~ inbuffer_data[608];
assign xnor5[609] = 1'b1 ^~ inbuffer_data[609];
assign xnor5[610] = 1'b1 ^~ inbuffer_data[610];
assign xnor5[611] = 1'b1 ^~ inbuffer_data[611];
assign xnor5[612] = 1'b0 ^~ inbuffer_data[612];
assign xnor5[613] = 1'b1 ^~ inbuffer_data[613];
assign xnor5[614] = 1'b1 ^~ inbuffer_data[614];
assign xnor5[615] = 1'b0 ^~ inbuffer_data[615];
assign xnor5[616] = 1'b0 ^~ inbuffer_data[616];
assign xnor5[617] = 1'b0 ^~ inbuffer_data[617];
assign xnor5[618] = 1'b1 ^~ inbuffer_data[618];
assign xnor5[619] = 1'b0 ^~ inbuffer_data[619];
assign xnor5[620] = 1'b1 ^~ inbuffer_data[620];
assign xnor5[621] = 1'b1 ^~ inbuffer_data[621];
assign xnor5[622] = 1'b0 ^~ inbuffer_data[622];
assign xnor5[623] = 1'b0 ^~ inbuffer_data[623];
assign xnor5[624] = 1'b1 ^~ inbuffer_data[624];
assign xnor5[625] = 1'b0 ^~ inbuffer_data[625];
assign xnor5[626] = 1'b1 ^~ inbuffer_data[626];
assign xnor5[627] = 1'b1 ^~ inbuffer_data[627];
assign xnor5[628] = 1'b1 ^~ inbuffer_data[628];
assign xnor5[629] = 1'b1 ^~ inbuffer_data[629];
assign xnor5[630] = 1'b1 ^~ inbuffer_data[630];
assign xnor5[631] = 1'b0 ^~ inbuffer_data[631];
assign xnor5[632] = 1'b1 ^~ inbuffer_data[632];
assign xnor5[633] = 1'b1 ^~ inbuffer_data[633];
assign xnor5[634] = 1'b1 ^~ inbuffer_data[634];
assign xnor5[635] = 1'b0 ^~ inbuffer_data[635];
assign xnor5[636] = 1'b1 ^~ inbuffer_data[636];
assign xnor5[637] = 1'b1 ^~ inbuffer_data[637];
assign xnor5[638] = 1'b1 ^~ inbuffer_data[638];
assign xnor5[639] = 1'b0 ^~ inbuffer_data[639];
assign xnor5[640] = 1'b1 ^~ inbuffer_data[640];
assign xnor5[641] = 1'b0 ^~ inbuffer_data[641];
assign xnor5[642] = 1'b0 ^~ inbuffer_data[642];
assign xnor5[643] = 1'b0 ^~ inbuffer_data[643];
assign xnor5[644] = 1'b1 ^~ inbuffer_data[644];
assign xnor5[645] = 1'b0 ^~ inbuffer_data[645];
assign xnor5[646] = 1'b1 ^~ inbuffer_data[646];
assign xnor5[647] = 1'b1 ^~ inbuffer_data[647];
assign xnor5[648] = 1'b1 ^~ inbuffer_data[648];
assign xnor5[649] = 1'b1 ^~ inbuffer_data[649];
assign xnor5[650] = 1'b0 ^~ inbuffer_data[650];
assign xnor5[651] = 1'b1 ^~ inbuffer_data[651];
assign xnor5[652] = 1'b1 ^~ inbuffer_data[652];
assign xnor5[653] = 1'b1 ^~ inbuffer_data[653];
assign xnor5[654] = 1'b1 ^~ inbuffer_data[654];
assign xnor5[655] = 1'b1 ^~ inbuffer_data[655];
assign xnor5[656] = 1'b0 ^~ inbuffer_data[656];
assign xnor5[657] = 1'b0 ^~ inbuffer_data[657];
assign xnor5[658] = 1'b0 ^~ inbuffer_data[658];
assign xnor5[659] = 1'b1 ^~ inbuffer_data[659];
assign xnor5[660] = 1'b1 ^~ inbuffer_data[660];
assign xnor5[661] = 1'b1 ^~ inbuffer_data[661];
assign xnor5[662] = 1'b0 ^~ inbuffer_data[662];
assign xnor5[663] = 1'b1 ^~ inbuffer_data[663];
assign xnor5[664] = 1'b1 ^~ inbuffer_data[664];
assign xnor5[665] = 1'b0 ^~ inbuffer_data[665];
assign xnor5[666] = 1'b1 ^~ inbuffer_data[666];
assign xnor5[667] = 1'b1 ^~ inbuffer_data[667];
assign xnor5[668] = 1'b0 ^~ inbuffer_data[668];
assign xnor5[669] = 1'b1 ^~ inbuffer_data[669];
assign xnor5[670] = 1'b1 ^~ inbuffer_data[670];
assign xnor5[671] = 1'b0 ^~ inbuffer_data[671];
assign xnor5[672] = 1'b1 ^~ inbuffer_data[672];
assign xnor5[673] = 1'b1 ^~ inbuffer_data[673];
assign xnor5[674] = 1'b0 ^~ inbuffer_data[674];
assign xnor5[675] = 1'b0 ^~ inbuffer_data[675];
assign xnor5[676] = 1'b0 ^~ inbuffer_data[676];
assign xnor5[677] = 1'b0 ^~ inbuffer_data[677];
assign xnor5[678] = 1'b0 ^~ inbuffer_data[678];
assign xnor5[679] = 1'b1 ^~ inbuffer_data[679];
assign xnor5[680] = 1'b1 ^~ inbuffer_data[680];
assign xnor5[681] = 1'b1 ^~ inbuffer_data[681];
assign xnor5[682] = 1'b1 ^~ inbuffer_data[682];
assign xnor5[683] = 1'b1 ^~ inbuffer_data[683];
assign xnor5[684] = 1'b1 ^~ inbuffer_data[684];
assign xnor5[685] = 1'b1 ^~ inbuffer_data[685];
assign xnor5[686] = 1'b1 ^~ inbuffer_data[686];
assign xnor5[687] = 1'b1 ^~ inbuffer_data[687];
assign xnor5[688] = 1'b0 ^~ inbuffer_data[688];
assign xnor5[689] = 1'b1 ^~ inbuffer_data[689];
assign xnor5[690] = 1'b0 ^~ inbuffer_data[690];
assign xnor5[691] = 1'b1 ^~ inbuffer_data[691];
assign xnor5[692] = 1'b0 ^~ inbuffer_data[692];
assign xnor5[693] = 1'b0 ^~ inbuffer_data[693];
assign xnor5[694] = 1'b0 ^~ inbuffer_data[694];
assign xnor5[695] = 1'b1 ^~ inbuffer_data[695];
assign xnor5[696] = 1'b0 ^~ inbuffer_data[696];
assign xnor5[697] = 1'b1 ^~ inbuffer_data[697];
assign xnor5[698] = 1'b0 ^~ inbuffer_data[698];
assign xnor5[699] = 1'b1 ^~ inbuffer_data[699];
assign xnor5[700] = 1'b0 ^~ inbuffer_data[700];
assign xnor5[701] = 1'b1 ^~ inbuffer_data[701];
assign xnor5[702] = 1'b0 ^~ inbuffer_data[702];
assign xnor5[703] = 1'b0 ^~ inbuffer_data[703];
assign xnor5[704] = 1'b1 ^~ inbuffer_data[704];
assign xnor5[705] = 1'b0 ^~ inbuffer_data[705];
assign xnor5[706] = 1'b0 ^~ inbuffer_data[706];
assign xnor5[707] = 1'b1 ^~ inbuffer_data[707];
assign xnor5[708] = 1'b0 ^~ inbuffer_data[708];
assign xnor5[709] = 1'b1 ^~ inbuffer_data[709];
assign xnor5[710] = 1'b1 ^~ inbuffer_data[710];
assign xnor5[711] = 1'b0 ^~ inbuffer_data[711];
assign xnor5[712] = 1'b1 ^~ inbuffer_data[712];
assign xnor5[713] = 1'b0 ^~ inbuffer_data[713];
assign xnor5[714] = 1'b1 ^~ inbuffer_data[714];
assign xnor5[715] = 1'b1 ^~ inbuffer_data[715];
assign xnor5[716] = 1'b0 ^~ inbuffer_data[716];
assign xnor5[717] = 1'b1 ^~ inbuffer_data[717];
assign xnor5[718] = 1'b1 ^~ inbuffer_data[718];
assign xnor5[719] = 1'b1 ^~ inbuffer_data[719];
assign xnor5[720] = 1'b0 ^~ inbuffer_data[720];
assign xnor5[721] = 1'b1 ^~ inbuffer_data[721];
assign xnor5[722] = 1'b0 ^~ inbuffer_data[722];
assign xnor5[723] = 1'b1 ^~ inbuffer_data[723];
assign xnor5[724] = 1'b1 ^~ inbuffer_data[724];
assign xnor5[725] = 1'b0 ^~ inbuffer_data[725];
assign xnor5[726] = 1'b1 ^~ inbuffer_data[726];
assign xnor5[727] = 1'b0 ^~ inbuffer_data[727];
assign xnor5[728] = 1'b0 ^~ inbuffer_data[728];
assign xnor5[729] = 1'b0 ^~ inbuffer_data[729];
assign xnor5[730] = 1'b0 ^~ inbuffer_data[730];
assign xnor5[731] = 1'b0 ^~ inbuffer_data[731];
assign xnor5[732] = 1'b0 ^~ inbuffer_data[732];
assign xnor5[733] = 1'b0 ^~ inbuffer_data[733];
assign xnor5[734] = 1'b0 ^~ inbuffer_data[734];
assign xnor5[735] = 1'b0 ^~ inbuffer_data[735];
assign xnor5[736] = 1'b0 ^~ inbuffer_data[736];
assign xnor5[737] = 1'b1 ^~ inbuffer_data[737];
assign xnor5[738] = 1'b1 ^~ inbuffer_data[738];
assign xnor5[739] = 1'b0 ^~ inbuffer_data[739];
assign xnor5[740] = 1'b0 ^~ inbuffer_data[740];
assign xnor5[741] = 1'b1 ^~ inbuffer_data[741];
assign xnor5[742] = 1'b0 ^~ inbuffer_data[742];
assign xnor5[743] = 1'b1 ^~ inbuffer_data[743];
assign xnor5[744] = 1'b1 ^~ inbuffer_data[744];
assign xnor5[745] = 1'b0 ^~ inbuffer_data[745];
assign xnor5[746] = 1'b0 ^~ inbuffer_data[746];
assign xnor5[747] = 1'b0 ^~ inbuffer_data[747];
assign xnor5[748] = 1'b1 ^~ inbuffer_data[748];
assign xnor5[749] = 1'b0 ^~ inbuffer_data[749];
assign xnor5[750] = 1'b1 ^~ inbuffer_data[750];
assign xnor5[751] = 1'b0 ^~ inbuffer_data[751];
assign xnor5[752] = 1'b0 ^~ inbuffer_data[752];
assign xnor5[753] = 1'b1 ^~ inbuffer_data[753];
assign xnor5[754] = 1'b0 ^~ inbuffer_data[754];
assign xnor5[755] = 1'b1 ^~ inbuffer_data[755];
assign xnor5[756] = 1'b1 ^~ inbuffer_data[756];
assign xnor5[757] = 1'b0 ^~ inbuffer_data[757];
assign xnor5[758] = 1'b0 ^~ inbuffer_data[758];
assign xnor5[759] = 1'b0 ^~ inbuffer_data[759];
assign xnor5[760] = 1'b0 ^~ inbuffer_data[760];
assign xnor5[761] = 1'b1 ^~ inbuffer_data[761];
assign xnor5[762] = 1'b0 ^~ inbuffer_data[762];
assign xnor5[763] = 1'b0 ^~ inbuffer_data[763];
assign xnor5[764] = 1'b0 ^~ inbuffer_data[764];
assign xnor5[765] = 1'b0 ^~ inbuffer_data[765];
assign xnor5[766] = 1'b1 ^~ inbuffer_data[766];
assign xnor5[767] = 1'b1 ^~ inbuffer_data[767];
assign xnor5[768] = 1'b0 ^~ inbuffer_data[768];
assign xnor5[769] = 1'b1 ^~ inbuffer_data[769];
assign xnor5[770] = 1'b1 ^~ inbuffer_data[770];
assign xnor5[771] = 1'b1 ^~ inbuffer_data[771];
assign xnor5[772] = 1'b1 ^~ inbuffer_data[772];
assign xnor5[773] = 1'b1 ^~ inbuffer_data[773];
assign xnor5[774] = 1'b1 ^~ inbuffer_data[774];
assign xnor5[775] = 1'b1 ^~ inbuffer_data[775];
assign xnor5[776] = 1'b0 ^~ inbuffer_data[776];
assign xnor5[777] = 1'b0 ^~ inbuffer_data[777];
assign xnor5[778] = 1'b0 ^~ inbuffer_data[778];
assign xnor5[779] = 1'b0 ^~ inbuffer_data[779];
assign xnor5[780] = 1'b1 ^~ inbuffer_data[780];
assign xnor5[781] = 1'b0 ^~ inbuffer_data[781];
assign xnor5[782] = 1'b1 ^~ inbuffer_data[782];
assign xnor5[783] = 1'b0 ^~ inbuffer_data[783];
assign xnor6[0] = 1'b0 ^~ inbuffer_data[0];
assign xnor6[1] = 1'b1 ^~ inbuffer_data[1];
assign xnor6[2] = 1'b0 ^~ inbuffer_data[2];
assign xnor6[3] = 1'b1 ^~ inbuffer_data[3];
assign xnor6[4] = 1'b1 ^~ inbuffer_data[4];
assign xnor6[5] = 1'b0 ^~ inbuffer_data[5];
assign xnor6[6] = 1'b1 ^~ inbuffer_data[6];
assign xnor6[7] = 1'b0 ^~ inbuffer_data[7];
assign xnor6[8] = 1'b0 ^~ inbuffer_data[8];
assign xnor6[9] = 1'b0 ^~ inbuffer_data[9];
assign xnor6[10] = 1'b0 ^~ inbuffer_data[10];
assign xnor6[11] = 1'b0 ^~ inbuffer_data[11];
assign xnor6[12] = 1'b1 ^~ inbuffer_data[12];
assign xnor6[13] = 1'b1 ^~ inbuffer_data[13];
assign xnor6[14] = 1'b1 ^~ inbuffer_data[14];
assign xnor6[15] = 1'b0 ^~ inbuffer_data[15];
assign xnor6[16] = 1'b1 ^~ inbuffer_data[16];
assign xnor6[17] = 1'b1 ^~ inbuffer_data[17];
assign xnor6[18] = 1'b1 ^~ inbuffer_data[18];
assign xnor6[19] = 1'b1 ^~ inbuffer_data[19];
assign xnor6[20] = 1'b1 ^~ inbuffer_data[20];
assign xnor6[21] = 1'b1 ^~ inbuffer_data[21];
assign xnor6[22] = 1'b1 ^~ inbuffer_data[22];
assign xnor6[23] = 1'b0 ^~ inbuffer_data[23];
assign xnor6[24] = 1'b0 ^~ inbuffer_data[24];
assign xnor6[25] = 1'b1 ^~ inbuffer_data[25];
assign xnor6[26] = 1'b0 ^~ inbuffer_data[26];
assign xnor6[27] = 1'b1 ^~ inbuffer_data[27];
assign xnor6[28] = 1'b1 ^~ inbuffer_data[28];
assign xnor6[29] = 1'b0 ^~ inbuffer_data[29];
assign xnor6[30] = 1'b0 ^~ inbuffer_data[30];
assign xnor6[31] = 1'b0 ^~ inbuffer_data[31];
assign xnor6[32] = 1'b0 ^~ inbuffer_data[32];
assign xnor6[33] = 1'b1 ^~ inbuffer_data[33];
assign xnor6[34] = 1'b1 ^~ inbuffer_data[34];
assign xnor6[35] = 1'b0 ^~ inbuffer_data[35];
assign xnor6[36] = 1'b0 ^~ inbuffer_data[36];
assign xnor6[37] = 1'b1 ^~ inbuffer_data[37];
assign xnor6[38] = 1'b1 ^~ inbuffer_data[38];
assign xnor6[39] = 1'b1 ^~ inbuffer_data[39];
assign xnor6[40] = 1'b1 ^~ inbuffer_data[40];
assign xnor6[41] = 1'b1 ^~ inbuffer_data[41];
assign xnor6[42] = 1'b1 ^~ inbuffer_data[42];
assign xnor6[43] = 1'b1 ^~ inbuffer_data[43];
assign xnor6[44] = 1'b1 ^~ inbuffer_data[44];
assign xnor6[45] = 1'b1 ^~ inbuffer_data[45];
assign xnor6[46] = 1'b1 ^~ inbuffer_data[46];
assign xnor6[47] = 1'b1 ^~ inbuffer_data[47];
assign xnor6[48] = 1'b1 ^~ inbuffer_data[48];
assign xnor6[49] = 1'b1 ^~ inbuffer_data[49];
assign xnor6[50] = 1'b0 ^~ inbuffer_data[50];
assign xnor6[51] = 1'b0 ^~ inbuffer_data[51];
assign xnor6[52] = 1'b1 ^~ inbuffer_data[52];
assign xnor6[53] = 1'b0 ^~ inbuffer_data[53];
assign xnor6[54] = 1'b0 ^~ inbuffer_data[54];
assign xnor6[55] = 1'b1 ^~ inbuffer_data[55];
assign xnor6[56] = 1'b0 ^~ inbuffer_data[56];
assign xnor6[57] = 1'b1 ^~ inbuffer_data[57];
assign xnor6[58] = 1'b0 ^~ inbuffer_data[58];
assign xnor6[59] = 1'b1 ^~ inbuffer_data[59];
assign xnor6[60] = 1'b1 ^~ inbuffer_data[60];
assign xnor6[61] = 1'b0 ^~ inbuffer_data[61];
assign xnor6[62] = 1'b0 ^~ inbuffer_data[62];
assign xnor6[63] = 1'b1 ^~ inbuffer_data[63];
assign xnor6[64] = 1'b0 ^~ inbuffer_data[64];
assign xnor6[65] = 1'b1 ^~ inbuffer_data[65];
assign xnor6[66] = 1'b1 ^~ inbuffer_data[66];
assign xnor6[67] = 1'b1 ^~ inbuffer_data[67];
assign xnor6[68] = 1'b1 ^~ inbuffer_data[68];
assign xnor6[69] = 1'b1 ^~ inbuffer_data[69];
assign xnor6[70] = 1'b1 ^~ inbuffer_data[70];
assign xnor6[71] = 1'b1 ^~ inbuffer_data[71];
assign xnor6[72] = 1'b1 ^~ inbuffer_data[72];
assign xnor6[73] = 1'b1 ^~ inbuffer_data[73];
assign xnor6[74] = 1'b1 ^~ inbuffer_data[74];
assign xnor6[75] = 1'b1 ^~ inbuffer_data[75];
assign xnor6[76] = 1'b1 ^~ inbuffer_data[76];
assign xnor6[77] = 1'b1 ^~ inbuffer_data[77];
assign xnor6[78] = 1'b1 ^~ inbuffer_data[78];
assign xnor6[79] = 1'b0 ^~ inbuffer_data[79];
assign xnor6[80] = 1'b1 ^~ inbuffer_data[80];
assign xnor6[81] = 1'b0 ^~ inbuffer_data[81];
assign xnor6[82] = 1'b1 ^~ inbuffer_data[82];
assign xnor6[83] = 1'b0 ^~ inbuffer_data[83];
assign xnor6[84] = 1'b1 ^~ inbuffer_data[84];
assign xnor6[85] = 1'b1 ^~ inbuffer_data[85];
assign xnor6[86] = 1'b1 ^~ inbuffer_data[86];
assign xnor6[87] = 1'b1 ^~ inbuffer_data[87];
assign xnor6[88] = 1'b0 ^~ inbuffer_data[88];
assign xnor6[89] = 1'b1 ^~ inbuffer_data[89];
assign xnor6[90] = 1'b0 ^~ inbuffer_data[90];
assign xnor6[91] = 1'b1 ^~ inbuffer_data[91];
assign xnor6[92] = 1'b0 ^~ inbuffer_data[92];
assign xnor6[93] = 1'b1 ^~ inbuffer_data[93];
assign xnor6[94] = 1'b1 ^~ inbuffer_data[94];
assign xnor6[95] = 1'b1 ^~ inbuffer_data[95];
assign xnor6[96] = 1'b1 ^~ inbuffer_data[96];
assign xnor6[97] = 1'b1 ^~ inbuffer_data[97];
assign xnor6[98] = 1'b1 ^~ inbuffer_data[98];
assign xnor6[99] = 1'b1 ^~ inbuffer_data[99];
assign xnor6[100] = 1'b1 ^~ inbuffer_data[100];
assign xnor6[101] = 1'b1 ^~ inbuffer_data[101];
assign xnor6[102] = 1'b1 ^~ inbuffer_data[102];
assign xnor6[103] = 1'b1 ^~ inbuffer_data[103];
assign xnor6[104] = 1'b1 ^~ inbuffer_data[104];
assign xnor6[105] = 1'b1 ^~ inbuffer_data[105];
assign xnor6[106] = 1'b1 ^~ inbuffer_data[106];
assign xnor6[107] = 1'b1 ^~ inbuffer_data[107];
assign xnor6[108] = 1'b1 ^~ inbuffer_data[108];
assign xnor6[109] = 1'b0 ^~ inbuffer_data[109];
assign xnor6[110] = 1'b0 ^~ inbuffer_data[110];
assign xnor6[111] = 1'b1 ^~ inbuffer_data[111];
assign xnor6[112] = 1'b0 ^~ inbuffer_data[112];
assign xnor6[113] = 1'b0 ^~ inbuffer_data[113];
assign xnor6[114] = 1'b0 ^~ inbuffer_data[114];
assign xnor6[115] = 1'b0 ^~ inbuffer_data[115];
assign xnor6[116] = 1'b1 ^~ inbuffer_data[116];
assign xnor6[117] = 1'b0 ^~ inbuffer_data[117];
assign xnor6[118] = 1'b0 ^~ inbuffer_data[118];
assign xnor6[119] = 1'b1 ^~ inbuffer_data[119];
assign xnor6[120] = 1'b1 ^~ inbuffer_data[120];
assign xnor6[121] = 1'b1 ^~ inbuffer_data[121];
assign xnor6[122] = 1'b0 ^~ inbuffer_data[122];
assign xnor6[123] = 1'b0 ^~ inbuffer_data[123];
assign xnor6[124] = 1'b0 ^~ inbuffer_data[124];
assign xnor6[125] = 1'b0 ^~ inbuffer_data[125];
assign xnor6[126] = 1'b0 ^~ inbuffer_data[126];
assign xnor6[127] = 1'b1 ^~ inbuffer_data[127];
assign xnor6[128] = 1'b1 ^~ inbuffer_data[128];
assign xnor6[129] = 1'b1 ^~ inbuffer_data[129];
assign xnor6[130] = 1'b1 ^~ inbuffer_data[130];
assign xnor6[131] = 1'b1 ^~ inbuffer_data[131];
assign xnor6[132] = 1'b1 ^~ inbuffer_data[132];
assign xnor6[133] = 1'b1 ^~ inbuffer_data[133];
assign xnor6[134] = 1'b1 ^~ inbuffer_data[134];
assign xnor6[135] = 1'b1 ^~ inbuffer_data[135];
assign xnor6[136] = 1'b0 ^~ inbuffer_data[136];
assign xnor6[137] = 1'b1 ^~ inbuffer_data[137];
assign xnor6[138] = 1'b1 ^~ inbuffer_data[138];
assign xnor6[139] = 1'b1 ^~ inbuffer_data[139];
assign xnor6[140] = 1'b1 ^~ inbuffer_data[140];
assign xnor6[141] = 1'b1 ^~ inbuffer_data[141];
assign xnor6[142] = 1'b1 ^~ inbuffer_data[142];
assign xnor6[143] = 1'b0 ^~ inbuffer_data[143];
assign xnor6[144] = 1'b1 ^~ inbuffer_data[144];
assign xnor6[145] = 1'b0 ^~ inbuffer_data[145];
assign xnor6[146] = 1'b1 ^~ inbuffer_data[146];
assign xnor6[147] = 1'b0 ^~ inbuffer_data[147];
assign xnor6[148] = 1'b1 ^~ inbuffer_data[148];
assign xnor6[149] = 1'b0 ^~ inbuffer_data[149];
assign xnor6[150] = 1'b1 ^~ inbuffer_data[150];
assign xnor6[151] = 1'b0 ^~ inbuffer_data[151];
assign xnor6[152] = 1'b0 ^~ inbuffer_data[152];
assign xnor6[153] = 1'b0 ^~ inbuffer_data[153];
assign xnor6[154] = 1'b1 ^~ inbuffer_data[154];
assign xnor6[155] = 1'b1 ^~ inbuffer_data[155];
assign xnor6[156] = 1'b0 ^~ inbuffer_data[156];
assign xnor6[157] = 1'b1 ^~ inbuffer_data[157];
assign xnor6[158] = 1'b1 ^~ inbuffer_data[158];
assign xnor6[159] = 1'b1 ^~ inbuffer_data[159];
assign xnor6[160] = 1'b1 ^~ inbuffer_data[160];
assign xnor6[161] = 1'b1 ^~ inbuffer_data[161];
assign xnor6[162] = 1'b1 ^~ inbuffer_data[162];
assign xnor6[163] = 1'b1 ^~ inbuffer_data[163];
assign xnor6[164] = 1'b1 ^~ inbuffer_data[164];
assign xnor6[165] = 1'b0 ^~ inbuffer_data[165];
assign xnor6[166] = 1'b1 ^~ inbuffer_data[166];
assign xnor6[167] = 1'b1 ^~ inbuffer_data[167];
assign xnor6[168] = 1'b0 ^~ inbuffer_data[168];
assign xnor6[169] = 1'b1 ^~ inbuffer_data[169];
assign xnor6[170] = 1'b0 ^~ inbuffer_data[170];
assign xnor6[171] = 1'b0 ^~ inbuffer_data[171];
assign xnor6[172] = 1'b1 ^~ inbuffer_data[172];
assign xnor6[173] = 1'b0 ^~ inbuffer_data[173];
assign xnor6[174] = 1'b1 ^~ inbuffer_data[174];
assign xnor6[175] = 1'b1 ^~ inbuffer_data[175];
assign xnor6[176] = 1'b0 ^~ inbuffer_data[176];
assign xnor6[177] = 1'b0 ^~ inbuffer_data[177];
assign xnor6[178] = 1'b0 ^~ inbuffer_data[178];
assign xnor6[179] = 1'b0 ^~ inbuffer_data[179];
assign xnor6[180] = 1'b0 ^~ inbuffer_data[180];
assign xnor6[181] = 1'b0 ^~ inbuffer_data[181];
assign xnor6[182] = 1'b0 ^~ inbuffer_data[182];
assign xnor6[183] = 1'b0 ^~ inbuffer_data[183];
assign xnor6[184] = 1'b1 ^~ inbuffer_data[184];
assign xnor6[185] = 1'b0 ^~ inbuffer_data[185];
assign xnor6[186] = 1'b0 ^~ inbuffer_data[186];
assign xnor6[187] = 1'b0 ^~ inbuffer_data[187];
assign xnor6[188] = 1'b1 ^~ inbuffer_data[188];
assign xnor6[189] = 1'b0 ^~ inbuffer_data[189];
assign xnor6[190] = 1'b0 ^~ inbuffer_data[190];
assign xnor6[191] = 1'b1 ^~ inbuffer_data[191];
assign xnor6[192] = 1'b0 ^~ inbuffer_data[192];
assign xnor6[193] = 1'b1 ^~ inbuffer_data[193];
assign xnor6[194] = 1'b0 ^~ inbuffer_data[194];
assign xnor6[195] = 1'b0 ^~ inbuffer_data[195];
assign xnor6[196] = 1'b0 ^~ inbuffer_data[196];
assign xnor6[197] = 1'b1 ^~ inbuffer_data[197];
assign xnor6[198] = 1'b0 ^~ inbuffer_data[198];
assign xnor6[199] = 1'b0 ^~ inbuffer_data[199];
assign xnor6[200] = 1'b1 ^~ inbuffer_data[200];
assign xnor6[201] = 1'b0 ^~ inbuffer_data[201];
assign xnor6[202] = 1'b0 ^~ inbuffer_data[202];
assign xnor6[203] = 1'b1 ^~ inbuffer_data[203];
assign xnor6[204] = 1'b0 ^~ inbuffer_data[204];
assign xnor6[205] = 1'b1 ^~ inbuffer_data[205];
assign xnor6[206] = 1'b1 ^~ inbuffer_data[206];
assign xnor6[207] = 1'b1 ^~ inbuffer_data[207];
assign xnor6[208] = 1'b0 ^~ inbuffer_data[208];
assign xnor6[209] = 1'b0 ^~ inbuffer_data[209];
assign xnor6[210] = 1'b0 ^~ inbuffer_data[210];
assign xnor6[211] = 1'b0 ^~ inbuffer_data[211];
assign xnor6[212] = 1'b0 ^~ inbuffer_data[212];
assign xnor6[213] = 1'b0 ^~ inbuffer_data[213];
assign xnor6[214] = 1'b0 ^~ inbuffer_data[214];
assign xnor6[215] = 1'b0 ^~ inbuffer_data[215];
assign xnor6[216] = 1'b0 ^~ inbuffer_data[216];
assign xnor6[217] = 1'b1 ^~ inbuffer_data[217];
assign xnor6[218] = 1'b0 ^~ inbuffer_data[218];
assign xnor6[219] = 1'b0 ^~ inbuffer_data[219];
assign xnor6[220] = 1'b1 ^~ inbuffer_data[220];
assign xnor6[221] = 1'b0 ^~ inbuffer_data[221];
assign xnor6[222] = 1'b0 ^~ inbuffer_data[222];
assign xnor6[223] = 1'b0 ^~ inbuffer_data[223];
assign xnor6[224] = 1'b0 ^~ inbuffer_data[224];
assign xnor6[225] = 1'b1 ^~ inbuffer_data[225];
assign xnor6[226] = 1'b0 ^~ inbuffer_data[226];
assign xnor6[227] = 1'b0 ^~ inbuffer_data[227];
assign xnor6[228] = 1'b0 ^~ inbuffer_data[228];
assign xnor6[229] = 1'b0 ^~ inbuffer_data[229];
assign xnor6[230] = 1'b0 ^~ inbuffer_data[230];
assign xnor6[231] = 1'b0 ^~ inbuffer_data[231];
assign xnor6[232] = 1'b0 ^~ inbuffer_data[232];
assign xnor6[233] = 1'b1 ^~ inbuffer_data[233];
assign xnor6[234] = 1'b1 ^~ inbuffer_data[234];
assign xnor6[235] = 1'b1 ^~ inbuffer_data[235];
assign xnor6[236] = 1'b1 ^~ inbuffer_data[236];
assign xnor6[237] = 1'b0 ^~ inbuffer_data[237];
assign xnor6[238] = 1'b0 ^~ inbuffer_data[238];
assign xnor6[239] = 1'b0 ^~ inbuffer_data[239];
assign xnor6[240] = 1'b0 ^~ inbuffer_data[240];
assign xnor6[241] = 1'b0 ^~ inbuffer_data[241];
assign xnor6[242] = 1'b0 ^~ inbuffer_data[242];
assign xnor6[243] = 1'b0 ^~ inbuffer_data[243];
assign xnor6[244] = 1'b0 ^~ inbuffer_data[244];
assign xnor6[245] = 1'b0 ^~ inbuffer_data[245];
assign xnor6[246] = 1'b0 ^~ inbuffer_data[246];
assign xnor6[247] = 1'b0 ^~ inbuffer_data[247];
assign xnor6[248] = 1'b0 ^~ inbuffer_data[248];
assign xnor6[249] = 1'b0 ^~ inbuffer_data[249];
assign xnor6[250] = 1'b0 ^~ inbuffer_data[250];
assign xnor6[251] = 1'b1 ^~ inbuffer_data[251];
assign xnor6[252] = 1'b0 ^~ inbuffer_data[252];
assign xnor6[253] = 1'b1 ^~ inbuffer_data[253];
assign xnor6[254] = 1'b1 ^~ inbuffer_data[254];
assign xnor6[255] = 1'b0 ^~ inbuffer_data[255];
assign xnor6[256] = 1'b0 ^~ inbuffer_data[256];
assign xnor6[257] = 1'b0 ^~ inbuffer_data[257];
assign xnor6[258] = 1'b0 ^~ inbuffer_data[258];
assign xnor6[259] = 1'b0 ^~ inbuffer_data[259];
assign xnor6[260] = 1'b1 ^~ inbuffer_data[260];
assign xnor6[261] = 1'b0 ^~ inbuffer_data[261];
assign xnor6[262] = 1'b0 ^~ inbuffer_data[262];
assign xnor6[263] = 1'b0 ^~ inbuffer_data[263];
assign xnor6[264] = 1'b0 ^~ inbuffer_data[264];
assign xnor6[265] = 1'b0 ^~ inbuffer_data[265];
assign xnor6[266] = 1'b0 ^~ inbuffer_data[266];
assign xnor6[267] = 1'b0 ^~ inbuffer_data[267];
assign xnor6[268] = 1'b0 ^~ inbuffer_data[268];
assign xnor6[269] = 1'b0 ^~ inbuffer_data[269];
assign xnor6[270] = 1'b0 ^~ inbuffer_data[270];
assign xnor6[271] = 1'b0 ^~ inbuffer_data[271];
assign xnor6[272] = 1'b0 ^~ inbuffer_data[272];
assign xnor6[273] = 1'b0 ^~ inbuffer_data[273];
assign xnor6[274] = 1'b0 ^~ inbuffer_data[274];
assign xnor6[275] = 1'b0 ^~ inbuffer_data[275];
assign xnor6[276] = 1'b0 ^~ inbuffer_data[276];
assign xnor6[277] = 1'b0 ^~ inbuffer_data[277];
assign xnor6[278] = 1'b0 ^~ inbuffer_data[278];
assign xnor6[279] = 1'b0 ^~ inbuffer_data[279];
assign xnor6[280] = 1'b1 ^~ inbuffer_data[280];
assign xnor6[281] = 1'b1 ^~ inbuffer_data[281];
assign xnor6[282] = 1'b1 ^~ inbuffer_data[282];
assign xnor6[283] = 1'b0 ^~ inbuffer_data[283];
assign xnor6[284] = 1'b0 ^~ inbuffer_data[284];
assign xnor6[285] = 1'b0 ^~ inbuffer_data[285];
assign xnor6[286] = 1'b0 ^~ inbuffer_data[286];
assign xnor6[287] = 1'b1 ^~ inbuffer_data[287];
assign xnor6[288] = 1'b0 ^~ inbuffer_data[288];
assign xnor6[289] = 1'b1 ^~ inbuffer_data[289];
assign xnor6[290] = 1'b0 ^~ inbuffer_data[290];
assign xnor6[291] = 1'b1 ^~ inbuffer_data[291];
assign xnor6[292] = 1'b0 ^~ inbuffer_data[292];
assign xnor6[293] = 1'b1 ^~ inbuffer_data[293];
assign xnor6[294] = 1'b0 ^~ inbuffer_data[294];
assign xnor6[295] = 1'b0 ^~ inbuffer_data[295];
assign xnor6[296] = 1'b0 ^~ inbuffer_data[296];
assign xnor6[297] = 1'b0 ^~ inbuffer_data[297];
assign xnor6[298] = 1'b0 ^~ inbuffer_data[298];
assign xnor6[299] = 1'b0 ^~ inbuffer_data[299];
assign xnor6[300] = 1'b0 ^~ inbuffer_data[300];
assign xnor6[301] = 1'b0 ^~ inbuffer_data[301];
assign xnor6[302] = 1'b0 ^~ inbuffer_data[302];
assign xnor6[303] = 1'b0 ^~ inbuffer_data[303];
assign xnor6[304] = 1'b0 ^~ inbuffer_data[304];
assign xnor6[305] = 1'b0 ^~ inbuffer_data[305];
assign xnor6[306] = 1'b0 ^~ inbuffer_data[306];
assign xnor6[307] = 1'b0 ^~ inbuffer_data[307];
assign xnor6[308] = 1'b0 ^~ inbuffer_data[308];
assign xnor6[309] = 1'b1 ^~ inbuffer_data[309];
assign xnor6[310] = 1'b0 ^~ inbuffer_data[310];
assign xnor6[311] = 1'b0 ^~ inbuffer_data[311];
assign xnor6[312] = 1'b1 ^~ inbuffer_data[312];
assign xnor6[313] = 1'b0 ^~ inbuffer_data[313];
assign xnor6[314] = 1'b0 ^~ inbuffer_data[314];
assign xnor6[315] = 1'b1 ^~ inbuffer_data[315];
assign xnor6[316] = 1'b1 ^~ inbuffer_data[316];
assign xnor6[317] = 1'b1 ^~ inbuffer_data[317];
assign xnor6[318] = 1'b1 ^~ inbuffer_data[318];
assign xnor6[319] = 1'b1 ^~ inbuffer_data[319];
assign xnor6[320] = 1'b1 ^~ inbuffer_data[320];
assign xnor6[321] = 1'b1 ^~ inbuffer_data[321];
assign xnor6[322] = 1'b0 ^~ inbuffer_data[322];
assign xnor6[323] = 1'b0 ^~ inbuffer_data[323];
assign xnor6[324] = 1'b0 ^~ inbuffer_data[324];
assign xnor6[325] = 1'b0 ^~ inbuffer_data[325];
assign xnor6[326] = 1'b0 ^~ inbuffer_data[326];
assign xnor6[327] = 1'b1 ^~ inbuffer_data[327];
assign xnor6[328] = 1'b1 ^~ inbuffer_data[328];
assign xnor6[329] = 1'b1 ^~ inbuffer_data[329];
assign xnor6[330] = 1'b0 ^~ inbuffer_data[330];
assign xnor6[331] = 1'b1 ^~ inbuffer_data[331];
assign xnor6[332] = 1'b1 ^~ inbuffer_data[332];
assign xnor6[333] = 1'b0 ^~ inbuffer_data[333];
assign xnor6[334] = 1'b0 ^~ inbuffer_data[334];
assign xnor6[335] = 1'b0 ^~ inbuffer_data[335];
assign xnor6[336] = 1'b1 ^~ inbuffer_data[336];
assign xnor6[337] = 1'b1 ^~ inbuffer_data[337];
assign xnor6[338] = 1'b0 ^~ inbuffer_data[338];
assign xnor6[339] = 1'b0 ^~ inbuffer_data[339];
assign xnor6[340] = 1'b0 ^~ inbuffer_data[340];
assign xnor6[341] = 1'b0 ^~ inbuffer_data[341];
assign xnor6[342] = 1'b1 ^~ inbuffer_data[342];
assign xnor6[343] = 1'b1 ^~ inbuffer_data[343];
assign xnor6[344] = 1'b1 ^~ inbuffer_data[344];
assign xnor6[345] = 1'b1 ^~ inbuffer_data[345];
assign xnor6[346] = 1'b0 ^~ inbuffer_data[346];
assign xnor6[347] = 1'b1 ^~ inbuffer_data[347];
assign xnor6[348] = 1'b1 ^~ inbuffer_data[348];
assign xnor6[349] = 1'b1 ^~ inbuffer_data[349];
assign xnor6[350] = 1'b0 ^~ inbuffer_data[350];
assign xnor6[351] = 1'b0 ^~ inbuffer_data[351];
assign xnor6[352] = 1'b0 ^~ inbuffer_data[352];
assign xnor6[353] = 1'b0 ^~ inbuffer_data[353];
assign xnor6[354] = 1'b0 ^~ inbuffer_data[354];
assign xnor6[355] = 1'b0 ^~ inbuffer_data[355];
assign xnor6[356] = 1'b0 ^~ inbuffer_data[356];
assign xnor6[357] = 1'b1 ^~ inbuffer_data[357];
assign xnor6[358] = 1'b1 ^~ inbuffer_data[358];
assign xnor6[359] = 1'b1 ^~ inbuffer_data[359];
assign xnor6[360] = 1'b1 ^~ inbuffer_data[360];
assign xnor6[361] = 1'b0 ^~ inbuffer_data[361];
assign xnor6[362] = 1'b0 ^~ inbuffer_data[362];
assign xnor6[363] = 1'b0 ^~ inbuffer_data[363];
assign xnor6[364] = 1'b0 ^~ inbuffer_data[364];
assign xnor6[365] = 1'b1 ^~ inbuffer_data[365];
assign xnor6[366] = 1'b0 ^~ inbuffer_data[366];
assign xnor6[367] = 1'b0 ^~ inbuffer_data[367];
assign xnor6[368] = 1'b0 ^~ inbuffer_data[368];
assign xnor6[369] = 1'b1 ^~ inbuffer_data[369];
assign xnor6[370] = 1'b1 ^~ inbuffer_data[370];
assign xnor6[371] = 1'b1 ^~ inbuffer_data[371];
assign xnor6[372] = 1'b0 ^~ inbuffer_data[372];
assign xnor6[373] = 1'b1 ^~ inbuffer_data[373];
assign xnor6[374] = 1'b1 ^~ inbuffer_data[374];
assign xnor6[375] = 1'b1 ^~ inbuffer_data[375];
assign xnor6[376] = 1'b1 ^~ inbuffer_data[376];
assign xnor6[377] = 1'b1 ^~ inbuffer_data[377];
assign xnor6[378] = 1'b0 ^~ inbuffer_data[378];
assign xnor6[379] = 1'b1 ^~ inbuffer_data[379];
assign xnor6[380] = 1'b1 ^~ inbuffer_data[380];
assign xnor6[381] = 1'b0 ^~ inbuffer_data[381];
assign xnor6[382] = 1'b0 ^~ inbuffer_data[382];
assign xnor6[383] = 1'b0 ^~ inbuffer_data[383];
assign xnor6[384] = 1'b0 ^~ inbuffer_data[384];
assign xnor6[385] = 1'b1 ^~ inbuffer_data[385];
assign xnor6[386] = 1'b1 ^~ inbuffer_data[386];
assign xnor6[387] = 1'b1 ^~ inbuffer_data[387];
assign xnor6[388] = 1'b1 ^~ inbuffer_data[388];
assign xnor6[389] = 1'b1 ^~ inbuffer_data[389];
assign xnor6[390] = 1'b0 ^~ inbuffer_data[390];
assign xnor6[391] = 1'b0 ^~ inbuffer_data[391];
assign xnor6[392] = 1'b1 ^~ inbuffer_data[392];
assign xnor6[393] = 1'b0 ^~ inbuffer_data[393];
assign xnor6[394] = 1'b0 ^~ inbuffer_data[394];
assign xnor6[395] = 1'b1 ^~ inbuffer_data[395];
assign xnor6[396] = 1'b0 ^~ inbuffer_data[396];
assign xnor6[397] = 1'b1 ^~ inbuffer_data[397];
assign xnor6[398] = 1'b1 ^~ inbuffer_data[398];
assign xnor6[399] = 1'b0 ^~ inbuffer_data[399];
assign xnor6[400] = 1'b1 ^~ inbuffer_data[400];
assign xnor6[401] = 1'b1 ^~ inbuffer_data[401];
assign xnor6[402] = 1'b1 ^~ inbuffer_data[402];
assign xnor6[403] = 1'b1 ^~ inbuffer_data[403];
assign xnor6[404] = 1'b1 ^~ inbuffer_data[404];
assign xnor6[405] = 1'b0 ^~ inbuffer_data[405];
assign xnor6[406] = 1'b0 ^~ inbuffer_data[406];
assign xnor6[407] = 1'b1 ^~ inbuffer_data[407];
assign xnor6[408] = 1'b1 ^~ inbuffer_data[408];
assign xnor6[409] = 1'b0 ^~ inbuffer_data[409];
assign xnor6[410] = 1'b1 ^~ inbuffer_data[410];
assign xnor6[411] = 1'b1 ^~ inbuffer_data[411];
assign xnor6[412] = 1'b1 ^~ inbuffer_data[412];
assign xnor6[413] = 1'b1 ^~ inbuffer_data[413];
assign xnor6[414] = 1'b1 ^~ inbuffer_data[414];
assign xnor6[415] = 1'b1 ^~ inbuffer_data[415];
assign xnor6[416] = 1'b1 ^~ inbuffer_data[416];
assign xnor6[417] = 1'b0 ^~ inbuffer_data[417];
assign xnor6[418] = 1'b1 ^~ inbuffer_data[418];
assign xnor6[419] = 1'b1 ^~ inbuffer_data[419];
assign xnor6[420] = 1'b0 ^~ inbuffer_data[420];
assign xnor6[421] = 1'b1 ^~ inbuffer_data[421];
assign xnor6[422] = 1'b1 ^~ inbuffer_data[422];
assign xnor6[423] = 1'b1 ^~ inbuffer_data[423];
assign xnor6[424] = 1'b0 ^~ inbuffer_data[424];
assign xnor6[425] = 1'b1 ^~ inbuffer_data[425];
assign xnor6[426] = 1'b1 ^~ inbuffer_data[426];
assign xnor6[427] = 1'b1 ^~ inbuffer_data[427];
assign xnor6[428] = 1'b1 ^~ inbuffer_data[428];
assign xnor6[429] = 1'b1 ^~ inbuffer_data[429];
assign xnor6[430] = 1'b1 ^~ inbuffer_data[430];
assign xnor6[431] = 1'b1 ^~ inbuffer_data[431];
assign xnor6[432] = 1'b1 ^~ inbuffer_data[432];
assign xnor6[433] = 1'b0 ^~ inbuffer_data[433];
assign xnor6[434] = 1'b1 ^~ inbuffer_data[434];
assign xnor6[435] = 1'b1 ^~ inbuffer_data[435];
assign xnor6[436] = 1'b0 ^~ inbuffer_data[436];
assign xnor6[437] = 1'b0 ^~ inbuffer_data[437];
assign xnor6[438] = 1'b0 ^~ inbuffer_data[438];
assign xnor6[439] = 1'b1 ^~ inbuffer_data[439];
assign xnor6[440] = 1'b0 ^~ inbuffer_data[440];
assign xnor6[441] = 1'b1 ^~ inbuffer_data[441];
assign xnor6[442] = 1'b1 ^~ inbuffer_data[442];
assign xnor6[443] = 1'b1 ^~ inbuffer_data[443];
assign xnor6[444] = 1'b1 ^~ inbuffer_data[444];
assign xnor6[445] = 1'b1 ^~ inbuffer_data[445];
assign xnor6[446] = 1'b0 ^~ inbuffer_data[446];
assign xnor6[447] = 1'b1 ^~ inbuffer_data[447];
assign xnor6[448] = 1'b0 ^~ inbuffer_data[448];
assign xnor6[449] = 1'b0 ^~ inbuffer_data[449];
assign xnor6[450] = 1'b0 ^~ inbuffer_data[450];
assign xnor6[451] = 1'b0 ^~ inbuffer_data[451];
assign xnor6[452] = 1'b0 ^~ inbuffer_data[452];
assign xnor6[453] = 1'b0 ^~ inbuffer_data[453];
assign xnor6[454] = 1'b1 ^~ inbuffer_data[454];
assign xnor6[455] = 1'b1 ^~ inbuffer_data[455];
assign xnor6[456] = 1'b1 ^~ inbuffer_data[456];
assign xnor6[457] = 1'b1 ^~ inbuffer_data[457];
assign xnor6[458] = 1'b1 ^~ inbuffer_data[458];
assign xnor6[459] = 1'b1 ^~ inbuffer_data[459];
assign xnor6[460] = 1'b1 ^~ inbuffer_data[460];
assign xnor6[461] = 1'b1 ^~ inbuffer_data[461];
assign xnor6[462] = 1'b1 ^~ inbuffer_data[462];
assign xnor6[463] = 1'b1 ^~ inbuffer_data[463];
assign xnor6[464] = 1'b1 ^~ inbuffer_data[464];
assign xnor6[465] = 1'b1 ^~ inbuffer_data[465];
assign xnor6[466] = 1'b1 ^~ inbuffer_data[466];
assign xnor6[467] = 1'b1 ^~ inbuffer_data[467];
assign xnor6[468] = 1'b1 ^~ inbuffer_data[468];
assign xnor6[469] = 1'b1 ^~ inbuffer_data[469];
assign xnor6[470] = 1'b1 ^~ inbuffer_data[470];
assign xnor6[471] = 1'b1 ^~ inbuffer_data[471];
assign xnor6[472] = 1'b0 ^~ inbuffer_data[472];
assign xnor6[473] = 1'b0 ^~ inbuffer_data[473];
assign xnor6[474] = 1'b1 ^~ inbuffer_data[474];
assign xnor6[475] = 1'b0 ^~ inbuffer_data[475];
assign xnor6[476] = 1'b0 ^~ inbuffer_data[476];
assign xnor6[477] = 1'b1 ^~ inbuffer_data[477];
assign xnor6[478] = 1'b0 ^~ inbuffer_data[478];
assign xnor6[479] = 1'b1 ^~ inbuffer_data[479];
assign xnor6[480] = 1'b0 ^~ inbuffer_data[480];
assign xnor6[481] = 1'b0 ^~ inbuffer_data[481];
assign xnor6[482] = 1'b1 ^~ inbuffer_data[482];
assign xnor6[483] = 1'b1 ^~ inbuffer_data[483];
assign xnor6[484] = 1'b1 ^~ inbuffer_data[484];
assign xnor6[485] = 1'b1 ^~ inbuffer_data[485];
assign xnor6[486] = 1'b1 ^~ inbuffer_data[486];
assign xnor6[487] = 1'b1 ^~ inbuffer_data[487];
assign xnor6[488] = 1'b1 ^~ inbuffer_data[488];
assign xnor6[489] = 1'b1 ^~ inbuffer_data[489];
assign xnor6[490] = 1'b0 ^~ inbuffer_data[490];
assign xnor6[491] = 1'b0 ^~ inbuffer_data[491];
assign xnor6[492] = 1'b0 ^~ inbuffer_data[492];
assign xnor6[493] = 1'b1 ^~ inbuffer_data[493];
assign xnor6[494] = 1'b0 ^~ inbuffer_data[494];
assign xnor6[495] = 1'b1 ^~ inbuffer_data[495];
assign xnor6[496] = 1'b1 ^~ inbuffer_data[496];
assign xnor6[497] = 1'b0 ^~ inbuffer_data[497];
assign xnor6[498] = 1'b1 ^~ inbuffer_data[498];
assign xnor6[499] = 1'b0 ^~ inbuffer_data[499];
assign xnor6[500] = 1'b0 ^~ inbuffer_data[500];
assign xnor6[501] = 1'b0 ^~ inbuffer_data[501];
assign xnor6[502] = 1'b1 ^~ inbuffer_data[502];
assign xnor6[503] = 1'b0 ^~ inbuffer_data[503];
assign xnor6[504] = 1'b0 ^~ inbuffer_data[504];
assign xnor6[505] = 1'b1 ^~ inbuffer_data[505];
assign xnor6[506] = 1'b0 ^~ inbuffer_data[506];
assign xnor6[507] = 1'b0 ^~ inbuffer_data[507];
assign xnor6[508] = 1'b0 ^~ inbuffer_data[508];
assign xnor6[509] = 1'b0 ^~ inbuffer_data[509];
assign xnor6[510] = 1'b0 ^~ inbuffer_data[510];
assign xnor6[511] = 1'b1 ^~ inbuffer_data[511];
assign xnor6[512] = 1'b1 ^~ inbuffer_data[512];
assign xnor6[513] = 1'b1 ^~ inbuffer_data[513];
assign xnor6[514] = 1'b1 ^~ inbuffer_data[514];
assign xnor6[515] = 1'b1 ^~ inbuffer_data[515];
assign xnor6[516] = 1'b1 ^~ inbuffer_data[516];
assign xnor6[517] = 1'b1 ^~ inbuffer_data[517];
assign xnor6[518] = 1'b1 ^~ inbuffer_data[518];
assign xnor6[519] = 1'b1 ^~ inbuffer_data[519];
assign xnor6[520] = 1'b1 ^~ inbuffer_data[520];
assign xnor6[521] = 1'b1 ^~ inbuffer_data[521];
assign xnor6[522] = 1'b1 ^~ inbuffer_data[522];
assign xnor6[523] = 1'b0 ^~ inbuffer_data[523];
assign xnor6[524] = 1'b0 ^~ inbuffer_data[524];
assign xnor6[525] = 1'b1 ^~ inbuffer_data[525];
assign xnor6[526] = 1'b0 ^~ inbuffer_data[526];
assign xnor6[527] = 1'b1 ^~ inbuffer_data[527];
assign xnor6[528] = 1'b1 ^~ inbuffer_data[528];
assign xnor6[529] = 1'b0 ^~ inbuffer_data[529];
assign xnor6[530] = 1'b1 ^~ inbuffer_data[530];
assign xnor6[531] = 1'b0 ^~ inbuffer_data[531];
assign xnor6[532] = 1'b1 ^~ inbuffer_data[532];
assign xnor6[533] = 1'b0 ^~ inbuffer_data[533];
assign xnor6[534] = 1'b1 ^~ inbuffer_data[534];
assign xnor6[535] = 1'b0 ^~ inbuffer_data[535];
assign xnor6[536] = 1'b0 ^~ inbuffer_data[536];
assign xnor6[537] = 1'b0 ^~ inbuffer_data[537];
assign xnor6[538] = 1'b1 ^~ inbuffer_data[538];
assign xnor6[539] = 1'b1 ^~ inbuffer_data[539];
assign xnor6[540] = 1'b0 ^~ inbuffer_data[540];
assign xnor6[541] = 1'b1 ^~ inbuffer_data[541];
assign xnor6[542] = 1'b1 ^~ inbuffer_data[542];
assign xnor6[543] = 1'b1 ^~ inbuffer_data[543];
assign xnor6[544] = 1'b1 ^~ inbuffer_data[544];
assign xnor6[545] = 1'b1 ^~ inbuffer_data[545];
assign xnor6[546] = 1'b1 ^~ inbuffer_data[546];
assign xnor6[547] = 1'b0 ^~ inbuffer_data[547];
assign xnor6[548] = 1'b1 ^~ inbuffer_data[548];
assign xnor6[549] = 1'b1 ^~ inbuffer_data[549];
assign xnor6[550] = 1'b1 ^~ inbuffer_data[550];
assign xnor6[551] = 1'b0 ^~ inbuffer_data[551];
assign xnor6[552] = 1'b1 ^~ inbuffer_data[552];
assign xnor6[553] = 1'b1 ^~ inbuffer_data[553];
assign xnor6[554] = 1'b1 ^~ inbuffer_data[554];
assign xnor6[555] = 1'b0 ^~ inbuffer_data[555];
assign xnor6[556] = 1'b0 ^~ inbuffer_data[556];
assign xnor6[557] = 1'b0 ^~ inbuffer_data[557];
assign xnor6[558] = 1'b1 ^~ inbuffer_data[558];
assign xnor6[559] = 1'b0 ^~ inbuffer_data[559];
assign xnor6[560] = 1'b0 ^~ inbuffer_data[560];
assign xnor6[561] = 1'b0 ^~ inbuffer_data[561];
assign xnor6[562] = 1'b0 ^~ inbuffer_data[562];
assign xnor6[563] = 1'b1 ^~ inbuffer_data[563];
assign xnor6[564] = 1'b0 ^~ inbuffer_data[564];
assign xnor6[565] = 1'b0 ^~ inbuffer_data[565];
assign xnor6[566] = 1'b0 ^~ inbuffer_data[566];
assign xnor6[567] = 1'b0 ^~ inbuffer_data[567];
assign xnor6[568] = 1'b0 ^~ inbuffer_data[568];
assign xnor6[569] = 1'b1 ^~ inbuffer_data[569];
assign xnor6[570] = 1'b1 ^~ inbuffer_data[570];
assign xnor6[571] = 1'b1 ^~ inbuffer_data[571];
assign xnor6[572] = 1'b1 ^~ inbuffer_data[572];
assign xnor6[573] = 1'b1 ^~ inbuffer_data[573];
assign xnor6[574] = 1'b1 ^~ inbuffer_data[574];
assign xnor6[575] = 1'b1 ^~ inbuffer_data[575];
assign xnor6[576] = 1'b1 ^~ inbuffer_data[576];
assign xnor6[577] = 1'b1 ^~ inbuffer_data[577];
assign xnor6[578] = 1'b1 ^~ inbuffer_data[578];
assign xnor6[579] = 1'b1 ^~ inbuffer_data[579];
assign xnor6[580] = 1'b1 ^~ inbuffer_data[580];
assign xnor6[581] = 1'b0 ^~ inbuffer_data[581];
assign xnor6[582] = 1'b0 ^~ inbuffer_data[582];
assign xnor6[583] = 1'b1 ^~ inbuffer_data[583];
assign xnor6[584] = 1'b0 ^~ inbuffer_data[584];
assign xnor6[585] = 1'b0 ^~ inbuffer_data[585];
assign xnor6[586] = 1'b1 ^~ inbuffer_data[586];
assign xnor6[587] = 1'b1 ^~ inbuffer_data[587];
assign xnor6[588] = 1'b1 ^~ inbuffer_data[588];
assign xnor6[589] = 1'b0 ^~ inbuffer_data[589];
assign xnor6[590] = 1'b1 ^~ inbuffer_data[590];
assign xnor6[591] = 1'b1 ^~ inbuffer_data[591];
assign xnor6[592] = 1'b0 ^~ inbuffer_data[592];
assign xnor6[593] = 1'b0 ^~ inbuffer_data[593];
assign xnor6[594] = 1'b0 ^~ inbuffer_data[594];
assign xnor6[595] = 1'b1 ^~ inbuffer_data[595];
assign xnor6[596] = 1'b1 ^~ inbuffer_data[596];
assign xnor6[597] = 1'b0 ^~ inbuffer_data[597];
assign xnor6[598] = 1'b1 ^~ inbuffer_data[598];
assign xnor6[599] = 1'b1 ^~ inbuffer_data[599];
assign xnor6[600] = 1'b1 ^~ inbuffer_data[600];
assign xnor6[601] = 1'b1 ^~ inbuffer_data[601];
assign xnor6[602] = 1'b1 ^~ inbuffer_data[602];
assign xnor6[603] = 1'b1 ^~ inbuffer_data[603];
assign xnor6[604] = 1'b1 ^~ inbuffer_data[604];
assign xnor6[605] = 1'b1 ^~ inbuffer_data[605];
assign xnor6[606] = 1'b1 ^~ inbuffer_data[606];
assign xnor6[607] = 1'b1 ^~ inbuffer_data[607];
assign xnor6[608] = 1'b1 ^~ inbuffer_data[608];
assign xnor6[609] = 1'b0 ^~ inbuffer_data[609];
assign xnor6[610] = 1'b1 ^~ inbuffer_data[610];
assign xnor6[611] = 1'b0 ^~ inbuffer_data[611];
assign xnor6[612] = 1'b1 ^~ inbuffer_data[612];
assign xnor6[613] = 1'b1 ^~ inbuffer_data[613];
assign xnor6[614] = 1'b1 ^~ inbuffer_data[614];
assign xnor6[615] = 1'b0 ^~ inbuffer_data[615];
assign xnor6[616] = 1'b0 ^~ inbuffer_data[616];
assign xnor6[617] = 1'b1 ^~ inbuffer_data[617];
assign xnor6[618] = 1'b0 ^~ inbuffer_data[618];
assign xnor6[619] = 1'b1 ^~ inbuffer_data[619];
assign xnor6[620] = 1'b0 ^~ inbuffer_data[620];
assign xnor6[621] = 1'b0 ^~ inbuffer_data[621];
assign xnor6[622] = 1'b0 ^~ inbuffer_data[622];
assign xnor6[623] = 1'b0 ^~ inbuffer_data[623];
assign xnor6[624] = 1'b0 ^~ inbuffer_data[624];
assign xnor6[625] = 1'b0 ^~ inbuffer_data[625];
assign xnor6[626] = 1'b1 ^~ inbuffer_data[626];
assign xnor6[627] = 1'b0 ^~ inbuffer_data[627];
assign xnor6[628] = 1'b1 ^~ inbuffer_data[628];
assign xnor6[629] = 1'b1 ^~ inbuffer_data[629];
assign xnor6[630] = 1'b1 ^~ inbuffer_data[630];
assign xnor6[631] = 1'b1 ^~ inbuffer_data[631];
assign xnor6[632] = 1'b0 ^~ inbuffer_data[632];
assign xnor6[633] = 1'b1 ^~ inbuffer_data[633];
assign xnor6[634] = 1'b1 ^~ inbuffer_data[634];
assign xnor6[635] = 1'b0 ^~ inbuffer_data[635];
assign xnor6[636] = 1'b1 ^~ inbuffer_data[636];
assign xnor6[637] = 1'b1 ^~ inbuffer_data[637];
assign xnor6[638] = 1'b0 ^~ inbuffer_data[638];
assign xnor6[639] = 1'b0 ^~ inbuffer_data[639];
assign xnor6[640] = 1'b0 ^~ inbuffer_data[640];
assign xnor6[641] = 1'b0 ^~ inbuffer_data[641];
assign xnor6[642] = 1'b0 ^~ inbuffer_data[642];
assign xnor6[643] = 1'b0 ^~ inbuffer_data[643];
assign xnor6[644] = 1'b1 ^~ inbuffer_data[644];
assign xnor6[645] = 1'b1 ^~ inbuffer_data[645];
assign xnor6[646] = 1'b1 ^~ inbuffer_data[646];
assign xnor6[647] = 1'b1 ^~ inbuffer_data[647];
assign xnor6[648] = 1'b0 ^~ inbuffer_data[648];
assign xnor6[649] = 1'b0 ^~ inbuffer_data[649];
assign xnor6[650] = 1'b1 ^~ inbuffer_data[650];
assign xnor6[651] = 1'b0 ^~ inbuffer_data[651];
assign xnor6[652] = 1'b0 ^~ inbuffer_data[652];
assign xnor6[653] = 1'b0 ^~ inbuffer_data[653];
assign xnor6[654] = 1'b0 ^~ inbuffer_data[654];
assign xnor6[655] = 1'b0 ^~ inbuffer_data[655];
assign xnor6[656] = 1'b0 ^~ inbuffer_data[656];
assign xnor6[657] = 1'b0 ^~ inbuffer_data[657];
assign xnor6[658] = 1'b0 ^~ inbuffer_data[658];
assign xnor6[659] = 1'b0 ^~ inbuffer_data[659];
assign xnor6[660] = 1'b0 ^~ inbuffer_data[660];
assign xnor6[661] = 1'b0 ^~ inbuffer_data[661];
assign xnor6[662] = 1'b0 ^~ inbuffer_data[662];
assign xnor6[663] = 1'b0 ^~ inbuffer_data[663];
assign xnor6[664] = 1'b1 ^~ inbuffer_data[664];
assign xnor6[665] = 1'b0 ^~ inbuffer_data[665];
assign xnor6[666] = 1'b0 ^~ inbuffer_data[666];
assign xnor6[667] = 1'b0 ^~ inbuffer_data[667];
assign xnor6[668] = 1'b1 ^~ inbuffer_data[668];
assign xnor6[669] = 1'b1 ^~ inbuffer_data[669];
assign xnor6[670] = 1'b0 ^~ inbuffer_data[670];
assign xnor6[671] = 1'b1 ^~ inbuffer_data[671];
assign xnor6[672] = 1'b1 ^~ inbuffer_data[672];
assign xnor6[673] = 1'b1 ^~ inbuffer_data[673];
assign xnor6[674] = 1'b0 ^~ inbuffer_data[674];
assign xnor6[675] = 1'b0 ^~ inbuffer_data[675];
assign xnor6[676] = 1'b0 ^~ inbuffer_data[676];
assign xnor6[677] = 1'b0 ^~ inbuffer_data[677];
assign xnor6[678] = 1'b0 ^~ inbuffer_data[678];
assign xnor6[679] = 1'b0 ^~ inbuffer_data[679];
assign xnor6[680] = 1'b0 ^~ inbuffer_data[680];
assign xnor6[681] = 1'b0 ^~ inbuffer_data[681];
assign xnor6[682] = 1'b0 ^~ inbuffer_data[682];
assign xnor6[683] = 1'b0 ^~ inbuffer_data[683];
assign xnor6[684] = 1'b0 ^~ inbuffer_data[684];
assign xnor6[685] = 1'b0 ^~ inbuffer_data[685];
assign xnor6[686] = 1'b0 ^~ inbuffer_data[686];
assign xnor6[687] = 1'b0 ^~ inbuffer_data[687];
assign xnor6[688] = 1'b0 ^~ inbuffer_data[688];
assign xnor6[689] = 1'b1 ^~ inbuffer_data[689];
assign xnor6[690] = 1'b0 ^~ inbuffer_data[690];
assign xnor6[691] = 1'b1 ^~ inbuffer_data[691];
assign xnor6[692] = 1'b0 ^~ inbuffer_data[692];
assign xnor6[693] = 1'b1 ^~ inbuffer_data[693];
assign xnor6[694] = 1'b0 ^~ inbuffer_data[694];
assign xnor6[695] = 1'b1 ^~ inbuffer_data[695];
assign xnor6[696] = 1'b1 ^~ inbuffer_data[696];
assign xnor6[697] = 1'b1 ^~ inbuffer_data[697];
assign xnor6[698] = 1'b1 ^~ inbuffer_data[698];
assign xnor6[699] = 1'b0 ^~ inbuffer_data[699];
assign xnor6[700] = 1'b1 ^~ inbuffer_data[700];
assign xnor6[701] = 1'b1 ^~ inbuffer_data[701];
assign xnor6[702] = 1'b0 ^~ inbuffer_data[702];
assign xnor6[703] = 1'b1 ^~ inbuffer_data[703];
assign xnor6[704] = 1'b0 ^~ inbuffer_data[704];
assign xnor6[705] = 1'b0 ^~ inbuffer_data[705];
assign xnor6[706] = 1'b0 ^~ inbuffer_data[706];
assign xnor6[707] = 1'b0 ^~ inbuffer_data[707];
assign xnor6[708] = 1'b0 ^~ inbuffer_data[708];
assign xnor6[709] = 1'b0 ^~ inbuffer_data[709];
assign xnor6[710] = 1'b1 ^~ inbuffer_data[710];
assign xnor6[711] = 1'b1 ^~ inbuffer_data[711];
assign xnor6[712] = 1'b0 ^~ inbuffer_data[712];
assign xnor6[713] = 1'b0 ^~ inbuffer_data[713];
assign xnor6[714] = 1'b0 ^~ inbuffer_data[714];
assign xnor6[715] = 1'b1 ^~ inbuffer_data[715];
assign xnor6[716] = 1'b1 ^~ inbuffer_data[716];
assign xnor6[717] = 1'b0 ^~ inbuffer_data[717];
assign xnor6[718] = 1'b0 ^~ inbuffer_data[718];
assign xnor6[719] = 1'b0 ^~ inbuffer_data[719];
assign xnor6[720] = 1'b0 ^~ inbuffer_data[720];
assign xnor6[721] = 1'b0 ^~ inbuffer_data[721];
assign xnor6[722] = 1'b0 ^~ inbuffer_data[722];
assign xnor6[723] = 1'b0 ^~ inbuffer_data[723];
assign xnor6[724] = 1'b1 ^~ inbuffer_data[724];
assign xnor6[725] = 1'b1 ^~ inbuffer_data[725];
assign xnor6[726] = 1'b1 ^~ inbuffer_data[726];
assign xnor6[727] = 1'b1 ^~ inbuffer_data[727];
assign xnor6[728] = 1'b0 ^~ inbuffer_data[728];
assign xnor6[729] = 1'b0 ^~ inbuffer_data[729];
assign xnor6[730] = 1'b0 ^~ inbuffer_data[730];
assign xnor6[731] = 1'b1 ^~ inbuffer_data[731];
assign xnor6[732] = 1'b1 ^~ inbuffer_data[732];
assign xnor6[733] = 1'b1 ^~ inbuffer_data[733];
assign xnor6[734] = 1'b0 ^~ inbuffer_data[734];
assign xnor6[735] = 1'b0 ^~ inbuffer_data[735];
assign xnor6[736] = 1'b0 ^~ inbuffer_data[736];
assign xnor6[737] = 1'b0 ^~ inbuffer_data[737];
assign xnor6[738] = 1'b0 ^~ inbuffer_data[738];
assign xnor6[739] = 1'b0 ^~ inbuffer_data[739];
assign xnor6[740] = 1'b1 ^~ inbuffer_data[740];
assign xnor6[741] = 1'b1 ^~ inbuffer_data[741];
assign xnor6[742] = 1'b1 ^~ inbuffer_data[742];
assign xnor6[743] = 1'b0 ^~ inbuffer_data[743];
assign xnor6[744] = 1'b1 ^~ inbuffer_data[744];
assign xnor6[745] = 1'b0 ^~ inbuffer_data[745];
assign xnor6[746] = 1'b1 ^~ inbuffer_data[746];
assign xnor6[747] = 1'b1 ^~ inbuffer_data[747];
assign xnor6[748] = 1'b0 ^~ inbuffer_data[748];
assign xnor6[749] = 1'b1 ^~ inbuffer_data[749];
assign xnor6[750] = 1'b1 ^~ inbuffer_data[750];
assign xnor6[751] = 1'b1 ^~ inbuffer_data[751];
assign xnor6[752] = 1'b0 ^~ inbuffer_data[752];
assign xnor6[753] = 1'b0 ^~ inbuffer_data[753];
assign xnor6[754] = 1'b1 ^~ inbuffer_data[754];
assign xnor6[755] = 1'b0 ^~ inbuffer_data[755];
assign xnor6[756] = 1'b1 ^~ inbuffer_data[756];
assign xnor6[757] = 1'b0 ^~ inbuffer_data[757];
assign xnor6[758] = 1'b0 ^~ inbuffer_data[758];
assign xnor6[759] = 1'b0 ^~ inbuffer_data[759];
assign xnor6[760] = 1'b1 ^~ inbuffer_data[760];
assign xnor6[761] = 1'b1 ^~ inbuffer_data[761];
assign xnor6[762] = 1'b0 ^~ inbuffer_data[762];
assign xnor6[763] = 1'b1 ^~ inbuffer_data[763];
assign xnor6[764] = 1'b0 ^~ inbuffer_data[764];
assign xnor6[765] = 1'b0 ^~ inbuffer_data[765];
assign xnor6[766] = 1'b0 ^~ inbuffer_data[766];
assign xnor6[767] = 1'b0 ^~ inbuffer_data[767];
assign xnor6[768] = 1'b1 ^~ inbuffer_data[768];
assign xnor6[769] = 1'b1 ^~ inbuffer_data[769];
assign xnor6[770] = 1'b0 ^~ inbuffer_data[770];
assign xnor6[771] = 1'b0 ^~ inbuffer_data[771];
assign xnor6[772] = 1'b1 ^~ inbuffer_data[772];
assign xnor6[773] = 1'b0 ^~ inbuffer_data[773];
assign xnor6[774] = 1'b1 ^~ inbuffer_data[774];
assign xnor6[775] = 1'b0 ^~ inbuffer_data[775];
assign xnor6[776] = 1'b0 ^~ inbuffer_data[776];
assign xnor6[777] = 1'b1 ^~ inbuffer_data[777];
assign xnor6[778] = 1'b0 ^~ inbuffer_data[778];
assign xnor6[779] = 1'b1 ^~ inbuffer_data[779];
assign xnor6[780] = 1'b0 ^~ inbuffer_data[780];
assign xnor6[781] = 1'b0 ^~ inbuffer_data[781];
assign xnor6[782] = 1'b0 ^~ inbuffer_data[782];
assign xnor6[783] = 1'b0 ^~ inbuffer_data[783];
assign xnor7[0] = 1'b1 ^~ inbuffer_data[0];
assign xnor7[1] = 1'b1 ^~ inbuffer_data[1];
assign xnor7[2] = 1'b1 ^~ inbuffer_data[2];
assign xnor7[3] = 1'b1 ^~ inbuffer_data[3];
assign xnor7[4] = 1'b0 ^~ inbuffer_data[4];
assign xnor7[5] = 1'b1 ^~ inbuffer_data[5];
assign xnor7[6] = 1'b1 ^~ inbuffer_data[6];
assign xnor7[7] = 1'b0 ^~ inbuffer_data[7];
assign xnor7[8] = 1'b1 ^~ inbuffer_data[8];
assign xnor7[9] = 1'b1 ^~ inbuffer_data[9];
assign xnor7[10] = 1'b1 ^~ inbuffer_data[10];
assign xnor7[11] = 1'b0 ^~ inbuffer_data[11];
assign xnor7[12] = 1'b1 ^~ inbuffer_data[12];
assign xnor7[13] = 1'b1 ^~ inbuffer_data[13];
assign xnor7[14] = 1'b1 ^~ inbuffer_data[14];
assign xnor7[15] = 1'b0 ^~ inbuffer_data[15];
assign xnor7[16] = 1'b0 ^~ inbuffer_data[16];
assign xnor7[17] = 1'b0 ^~ inbuffer_data[17];
assign xnor7[18] = 1'b1 ^~ inbuffer_data[18];
assign xnor7[19] = 1'b1 ^~ inbuffer_data[19];
assign xnor7[20] = 1'b1 ^~ inbuffer_data[20];
assign xnor7[21] = 1'b1 ^~ inbuffer_data[21];
assign xnor7[22] = 1'b1 ^~ inbuffer_data[22];
assign xnor7[23] = 1'b0 ^~ inbuffer_data[23];
assign xnor7[24] = 1'b0 ^~ inbuffer_data[24];
assign xnor7[25] = 1'b0 ^~ inbuffer_data[25];
assign xnor7[26] = 1'b0 ^~ inbuffer_data[26];
assign xnor7[27] = 1'b0 ^~ inbuffer_data[27];
assign xnor7[28] = 1'b0 ^~ inbuffer_data[28];
assign xnor7[29] = 1'b1 ^~ inbuffer_data[29];
assign xnor7[30] = 1'b1 ^~ inbuffer_data[30];
assign xnor7[31] = 1'b0 ^~ inbuffer_data[31];
assign xnor7[32] = 1'b1 ^~ inbuffer_data[32];
assign xnor7[33] = 1'b1 ^~ inbuffer_data[33];
assign xnor7[34] = 1'b1 ^~ inbuffer_data[34];
assign xnor7[35] = 1'b1 ^~ inbuffer_data[35];
assign xnor7[36] = 1'b0 ^~ inbuffer_data[36];
assign xnor7[37] = 1'b0 ^~ inbuffer_data[37];
assign xnor7[38] = 1'b0 ^~ inbuffer_data[38];
assign xnor7[39] = 1'b1 ^~ inbuffer_data[39];
assign xnor7[40] = 1'b0 ^~ inbuffer_data[40];
assign xnor7[41] = 1'b0 ^~ inbuffer_data[41];
assign xnor7[42] = 1'b0 ^~ inbuffer_data[42];
assign xnor7[43] = 1'b1 ^~ inbuffer_data[43];
assign xnor7[44] = 1'b0 ^~ inbuffer_data[44];
assign xnor7[45] = 1'b1 ^~ inbuffer_data[45];
assign xnor7[46] = 1'b0 ^~ inbuffer_data[46];
assign xnor7[47] = 1'b1 ^~ inbuffer_data[47];
assign xnor7[48] = 1'b1 ^~ inbuffer_data[48];
assign xnor7[49] = 1'b0 ^~ inbuffer_data[49];
assign xnor7[50] = 1'b1 ^~ inbuffer_data[50];
assign xnor7[51] = 1'b0 ^~ inbuffer_data[51];
assign xnor7[52] = 1'b0 ^~ inbuffer_data[52];
assign xnor7[53] = 1'b1 ^~ inbuffer_data[53];
assign xnor7[54] = 1'b1 ^~ inbuffer_data[54];
assign xnor7[55] = 1'b0 ^~ inbuffer_data[55];
assign xnor7[56] = 1'b0 ^~ inbuffer_data[56];
assign xnor7[57] = 1'b1 ^~ inbuffer_data[57];
assign xnor7[58] = 1'b0 ^~ inbuffer_data[58];
assign xnor7[59] = 1'b1 ^~ inbuffer_data[59];
assign xnor7[60] = 1'b1 ^~ inbuffer_data[60];
assign xnor7[61] = 1'b1 ^~ inbuffer_data[61];
assign xnor7[62] = 1'b0 ^~ inbuffer_data[62];
assign xnor7[63] = 1'b0 ^~ inbuffer_data[63];
assign xnor7[64] = 1'b0 ^~ inbuffer_data[64];
assign xnor7[65] = 1'b0 ^~ inbuffer_data[65];
assign xnor7[66] = 1'b0 ^~ inbuffer_data[66];
assign xnor7[67] = 1'b1 ^~ inbuffer_data[67];
assign xnor7[68] = 1'b0 ^~ inbuffer_data[68];
assign xnor7[69] = 1'b0 ^~ inbuffer_data[69];
assign xnor7[70] = 1'b0 ^~ inbuffer_data[70];
assign xnor7[71] = 1'b0 ^~ inbuffer_data[71];
assign xnor7[72] = 1'b0 ^~ inbuffer_data[72];
assign xnor7[73] = 1'b1 ^~ inbuffer_data[73];
assign xnor7[74] = 1'b1 ^~ inbuffer_data[74];
assign xnor7[75] = 1'b0 ^~ inbuffer_data[75];
assign xnor7[76] = 1'b0 ^~ inbuffer_data[76];
assign xnor7[77] = 1'b1 ^~ inbuffer_data[77];
assign xnor7[78] = 1'b0 ^~ inbuffer_data[78];
assign xnor7[79] = 1'b0 ^~ inbuffer_data[79];
assign xnor7[80] = 1'b0 ^~ inbuffer_data[80];
assign xnor7[81] = 1'b1 ^~ inbuffer_data[81];
assign xnor7[82] = 1'b0 ^~ inbuffer_data[82];
assign xnor7[83] = 1'b0 ^~ inbuffer_data[83];
assign xnor7[84] = 1'b1 ^~ inbuffer_data[84];
assign xnor7[85] = 1'b0 ^~ inbuffer_data[85];
assign xnor7[86] = 1'b1 ^~ inbuffer_data[86];
assign xnor7[87] = 1'b0 ^~ inbuffer_data[87];
assign xnor7[88] = 1'b0 ^~ inbuffer_data[88];
assign xnor7[89] = 1'b0 ^~ inbuffer_data[89];
assign xnor7[90] = 1'b0 ^~ inbuffer_data[90];
assign xnor7[91] = 1'b1 ^~ inbuffer_data[91];
assign xnor7[92] = 1'b1 ^~ inbuffer_data[92];
assign xnor7[93] = 1'b0 ^~ inbuffer_data[93];
assign xnor7[94] = 1'b0 ^~ inbuffer_data[94];
assign xnor7[95] = 1'b1 ^~ inbuffer_data[95];
assign xnor7[96] = 1'b0 ^~ inbuffer_data[96];
assign xnor7[97] = 1'b0 ^~ inbuffer_data[97];
assign xnor7[98] = 1'b1 ^~ inbuffer_data[98];
assign xnor7[99] = 1'b0 ^~ inbuffer_data[99];
assign xnor7[100] = 1'b1 ^~ inbuffer_data[100];
assign xnor7[101] = 1'b0 ^~ inbuffer_data[101];
assign xnor7[102] = 1'b1 ^~ inbuffer_data[102];
assign xnor7[103] = 1'b0 ^~ inbuffer_data[103];
assign xnor7[104] = 1'b1 ^~ inbuffer_data[104];
assign xnor7[105] = 1'b0 ^~ inbuffer_data[105];
assign xnor7[106] = 1'b0 ^~ inbuffer_data[106];
assign xnor7[107] = 1'b1 ^~ inbuffer_data[107];
assign xnor7[108] = 1'b0 ^~ inbuffer_data[108];
assign xnor7[109] = 1'b1 ^~ inbuffer_data[109];
assign xnor7[110] = 1'b0 ^~ inbuffer_data[110];
assign xnor7[111] = 1'b1 ^~ inbuffer_data[111];
assign xnor7[112] = 1'b1 ^~ inbuffer_data[112];
assign xnor7[113] = 1'b1 ^~ inbuffer_data[113];
assign xnor7[114] = 1'b0 ^~ inbuffer_data[114];
assign xnor7[115] = 1'b1 ^~ inbuffer_data[115];
assign xnor7[116] = 1'b0 ^~ inbuffer_data[116];
assign xnor7[117] = 1'b1 ^~ inbuffer_data[117];
assign xnor7[118] = 1'b0 ^~ inbuffer_data[118];
assign xnor7[119] = 1'b0 ^~ inbuffer_data[119];
assign xnor7[120] = 1'b1 ^~ inbuffer_data[120];
assign xnor7[121] = 1'b1 ^~ inbuffer_data[121];
assign xnor7[122] = 1'b0 ^~ inbuffer_data[122];
assign xnor7[123] = 1'b0 ^~ inbuffer_data[123];
assign xnor7[124] = 1'b0 ^~ inbuffer_data[124];
assign xnor7[125] = 1'b0 ^~ inbuffer_data[125];
assign xnor7[126] = 1'b0 ^~ inbuffer_data[126];
assign xnor7[127] = 1'b0 ^~ inbuffer_data[127];
assign xnor7[128] = 1'b0 ^~ inbuffer_data[128];
assign xnor7[129] = 1'b0 ^~ inbuffer_data[129];
assign xnor7[130] = 1'b0 ^~ inbuffer_data[130];
assign xnor7[131] = 1'b1 ^~ inbuffer_data[131];
assign xnor7[132] = 1'b0 ^~ inbuffer_data[132];
assign xnor7[133] = 1'b1 ^~ inbuffer_data[133];
assign xnor7[134] = 1'b1 ^~ inbuffer_data[134];
assign xnor7[135] = 1'b1 ^~ inbuffer_data[135];
assign xnor7[136] = 1'b0 ^~ inbuffer_data[136];
assign xnor7[137] = 1'b0 ^~ inbuffer_data[137];
assign xnor7[138] = 1'b0 ^~ inbuffer_data[138];
assign xnor7[139] = 1'b1 ^~ inbuffer_data[139];
assign xnor7[140] = 1'b1 ^~ inbuffer_data[140];
assign xnor7[141] = 1'b1 ^~ inbuffer_data[141];
assign xnor7[142] = 1'b1 ^~ inbuffer_data[142];
assign xnor7[143] = 1'b1 ^~ inbuffer_data[143];
assign xnor7[144] = 1'b1 ^~ inbuffer_data[144];
assign xnor7[145] = 1'b1 ^~ inbuffer_data[145];
assign xnor7[146] = 1'b0 ^~ inbuffer_data[146];
assign xnor7[147] = 1'b1 ^~ inbuffer_data[147];
assign xnor7[148] = 1'b0 ^~ inbuffer_data[148];
assign xnor7[149] = 1'b1 ^~ inbuffer_data[149];
assign xnor7[150] = 1'b0 ^~ inbuffer_data[150];
assign xnor7[151] = 1'b0 ^~ inbuffer_data[151];
assign xnor7[152] = 1'b0 ^~ inbuffer_data[152];
assign xnor7[153] = 1'b0 ^~ inbuffer_data[153];
assign xnor7[154] = 1'b0 ^~ inbuffer_data[154];
assign xnor7[155] = 1'b0 ^~ inbuffer_data[155];
assign xnor7[156] = 1'b0 ^~ inbuffer_data[156];
assign xnor7[157] = 1'b0 ^~ inbuffer_data[157];
assign xnor7[158] = 1'b0 ^~ inbuffer_data[158];
assign xnor7[159] = 1'b0 ^~ inbuffer_data[159];
assign xnor7[160] = 1'b0 ^~ inbuffer_data[160];
assign xnor7[161] = 1'b0 ^~ inbuffer_data[161];
assign xnor7[162] = 1'b0 ^~ inbuffer_data[162];
assign xnor7[163] = 1'b1 ^~ inbuffer_data[163];
assign xnor7[164] = 1'b0 ^~ inbuffer_data[164];
assign xnor7[165] = 1'b1 ^~ inbuffer_data[165];
assign xnor7[166] = 1'b1 ^~ inbuffer_data[166];
assign xnor7[167] = 1'b0 ^~ inbuffer_data[167];
assign xnor7[168] = 1'b0 ^~ inbuffer_data[168];
assign xnor7[169] = 1'b0 ^~ inbuffer_data[169];
assign xnor7[170] = 1'b1 ^~ inbuffer_data[170];
assign xnor7[171] = 1'b0 ^~ inbuffer_data[171];
assign xnor7[172] = 1'b0 ^~ inbuffer_data[172];
assign xnor7[173] = 1'b1 ^~ inbuffer_data[173];
assign xnor7[174] = 1'b1 ^~ inbuffer_data[174];
assign xnor7[175] = 1'b1 ^~ inbuffer_data[175];
assign xnor7[176] = 1'b1 ^~ inbuffer_data[176];
assign xnor7[177] = 1'b1 ^~ inbuffer_data[177];
assign xnor7[178] = 1'b1 ^~ inbuffer_data[178];
assign xnor7[179] = 1'b1 ^~ inbuffer_data[179];
assign xnor7[180] = 1'b1 ^~ inbuffer_data[180];
assign xnor7[181] = 1'b1 ^~ inbuffer_data[181];
assign xnor7[182] = 1'b0 ^~ inbuffer_data[182];
assign xnor7[183] = 1'b1 ^~ inbuffer_data[183];
assign xnor7[184] = 1'b1 ^~ inbuffer_data[184];
assign xnor7[185] = 1'b1 ^~ inbuffer_data[185];
assign xnor7[186] = 1'b1 ^~ inbuffer_data[186];
assign xnor7[187] = 1'b0 ^~ inbuffer_data[187];
assign xnor7[188] = 1'b0 ^~ inbuffer_data[188];
assign xnor7[189] = 1'b0 ^~ inbuffer_data[189];
assign xnor7[190] = 1'b1 ^~ inbuffer_data[190];
assign xnor7[191] = 1'b0 ^~ inbuffer_data[191];
assign xnor7[192] = 1'b0 ^~ inbuffer_data[192];
assign xnor7[193] = 1'b0 ^~ inbuffer_data[193];
assign xnor7[194] = 1'b0 ^~ inbuffer_data[194];
assign xnor7[195] = 1'b0 ^~ inbuffer_data[195];
assign xnor7[196] = 1'b0 ^~ inbuffer_data[196];
assign xnor7[197] = 1'b0 ^~ inbuffer_data[197];
assign xnor7[198] = 1'b0 ^~ inbuffer_data[198];
assign xnor7[199] = 1'b1 ^~ inbuffer_data[199];
assign xnor7[200] = 1'b1 ^~ inbuffer_data[200];
assign xnor7[201] = 1'b1 ^~ inbuffer_data[201];
assign xnor7[202] = 1'b1 ^~ inbuffer_data[202];
assign xnor7[203] = 1'b1 ^~ inbuffer_data[203];
assign xnor7[204] = 1'b1 ^~ inbuffer_data[204];
assign xnor7[205] = 1'b1 ^~ inbuffer_data[205];
assign xnor7[206] = 1'b1 ^~ inbuffer_data[206];
assign xnor7[207] = 1'b1 ^~ inbuffer_data[207];
assign xnor7[208] = 1'b1 ^~ inbuffer_data[208];
assign xnor7[209] = 1'b1 ^~ inbuffer_data[209];
assign xnor7[210] = 1'b0 ^~ inbuffer_data[210];
assign xnor7[211] = 1'b0 ^~ inbuffer_data[211];
assign xnor7[212] = 1'b0 ^~ inbuffer_data[212];
assign xnor7[213] = 1'b1 ^~ inbuffer_data[213];
assign xnor7[214] = 1'b1 ^~ inbuffer_data[214];
assign xnor7[215] = 1'b1 ^~ inbuffer_data[215];
assign xnor7[216] = 1'b1 ^~ inbuffer_data[216];
assign xnor7[217] = 1'b1 ^~ inbuffer_data[217];
assign xnor7[218] = 1'b0 ^~ inbuffer_data[218];
assign xnor7[219] = 1'b0 ^~ inbuffer_data[219];
assign xnor7[220] = 1'b0 ^~ inbuffer_data[220];
assign xnor7[221] = 1'b0 ^~ inbuffer_data[221];
assign xnor7[222] = 1'b1 ^~ inbuffer_data[222];
assign xnor7[223] = 1'b0 ^~ inbuffer_data[223];
assign xnor7[224] = 1'b1 ^~ inbuffer_data[224];
assign xnor7[225] = 1'b1 ^~ inbuffer_data[225];
assign xnor7[226] = 1'b0 ^~ inbuffer_data[226];
assign xnor7[227] = 1'b1 ^~ inbuffer_data[227];
assign xnor7[228] = 1'b1 ^~ inbuffer_data[228];
assign xnor7[229] = 1'b1 ^~ inbuffer_data[229];
assign xnor7[230] = 1'b1 ^~ inbuffer_data[230];
assign xnor7[231] = 1'b1 ^~ inbuffer_data[231];
assign xnor7[232] = 1'b1 ^~ inbuffer_data[232];
assign xnor7[233] = 1'b0 ^~ inbuffer_data[233];
assign xnor7[234] = 1'b1 ^~ inbuffer_data[234];
assign xnor7[235] = 1'b1 ^~ inbuffer_data[235];
assign xnor7[236] = 1'b1 ^~ inbuffer_data[236];
assign xnor7[237] = 1'b1 ^~ inbuffer_data[237];
assign xnor7[238] = 1'b1 ^~ inbuffer_data[238];
assign xnor7[239] = 1'b1 ^~ inbuffer_data[239];
assign xnor7[240] = 1'b1 ^~ inbuffer_data[240];
assign xnor7[241] = 1'b1 ^~ inbuffer_data[241];
assign xnor7[242] = 1'b1 ^~ inbuffer_data[242];
assign xnor7[243] = 1'b1 ^~ inbuffer_data[243];
assign xnor7[244] = 1'b1 ^~ inbuffer_data[244];
assign xnor7[245] = 1'b0 ^~ inbuffer_data[245];
assign xnor7[246] = 1'b1 ^~ inbuffer_data[246];
assign xnor7[247] = 1'b0 ^~ inbuffer_data[247];
assign xnor7[248] = 1'b0 ^~ inbuffer_data[248];
assign xnor7[249] = 1'b1 ^~ inbuffer_data[249];
assign xnor7[250] = 1'b0 ^~ inbuffer_data[250];
assign xnor7[251] = 1'b0 ^~ inbuffer_data[251];
assign xnor7[252] = 1'b0 ^~ inbuffer_data[252];
assign xnor7[253] = 1'b1 ^~ inbuffer_data[253];
assign xnor7[254] = 1'b1 ^~ inbuffer_data[254];
assign xnor7[255] = 1'b1 ^~ inbuffer_data[255];
assign xnor7[256] = 1'b1 ^~ inbuffer_data[256];
assign xnor7[257] = 1'b1 ^~ inbuffer_data[257];
assign xnor7[258] = 1'b1 ^~ inbuffer_data[258];
assign xnor7[259] = 1'b1 ^~ inbuffer_data[259];
assign xnor7[260] = 1'b1 ^~ inbuffer_data[260];
assign xnor7[261] = 1'b1 ^~ inbuffer_data[261];
assign xnor7[262] = 1'b0 ^~ inbuffer_data[262];
assign xnor7[263] = 1'b1 ^~ inbuffer_data[263];
assign xnor7[264] = 1'b1 ^~ inbuffer_data[264];
assign xnor7[265] = 1'b1 ^~ inbuffer_data[265];
assign xnor7[266] = 1'b1 ^~ inbuffer_data[266];
assign xnor7[267] = 1'b1 ^~ inbuffer_data[267];
assign xnor7[268] = 1'b1 ^~ inbuffer_data[268];
assign xnor7[269] = 1'b1 ^~ inbuffer_data[269];
assign xnor7[270] = 1'b1 ^~ inbuffer_data[270];
assign xnor7[271] = 1'b1 ^~ inbuffer_data[271];
assign xnor7[272] = 1'b1 ^~ inbuffer_data[272];
assign xnor7[273] = 1'b0 ^~ inbuffer_data[273];
assign xnor7[274] = 1'b0 ^~ inbuffer_data[274];
assign xnor7[275] = 1'b0 ^~ inbuffer_data[275];
assign xnor7[276] = 1'b0 ^~ inbuffer_data[276];
assign xnor7[277] = 1'b1 ^~ inbuffer_data[277];
assign xnor7[278] = 1'b0 ^~ inbuffer_data[278];
assign xnor7[279] = 1'b1 ^~ inbuffer_data[279];
assign xnor7[280] = 1'b0 ^~ inbuffer_data[280];
assign xnor7[281] = 1'b1 ^~ inbuffer_data[281];
assign xnor7[282] = 1'b1 ^~ inbuffer_data[282];
assign xnor7[283] = 1'b1 ^~ inbuffer_data[283];
assign xnor7[284] = 1'b1 ^~ inbuffer_data[284];
assign xnor7[285] = 1'b1 ^~ inbuffer_data[285];
assign xnor7[286] = 1'b1 ^~ inbuffer_data[286];
assign xnor7[287] = 1'b1 ^~ inbuffer_data[287];
assign xnor7[288] = 1'b1 ^~ inbuffer_data[288];
assign xnor7[289] = 1'b1 ^~ inbuffer_data[289];
assign xnor7[290] = 1'b1 ^~ inbuffer_data[290];
assign xnor7[291] = 1'b1 ^~ inbuffer_data[291];
assign xnor7[292] = 1'b1 ^~ inbuffer_data[292];
assign xnor7[293] = 1'b1 ^~ inbuffer_data[293];
assign xnor7[294] = 1'b1 ^~ inbuffer_data[294];
assign xnor7[295] = 1'b1 ^~ inbuffer_data[295];
assign xnor7[296] = 1'b1 ^~ inbuffer_data[296];
assign xnor7[297] = 1'b1 ^~ inbuffer_data[297];
assign xnor7[298] = 1'b1 ^~ inbuffer_data[298];
assign xnor7[299] = 1'b1 ^~ inbuffer_data[299];
assign xnor7[300] = 1'b1 ^~ inbuffer_data[300];
assign xnor7[301] = 1'b1 ^~ inbuffer_data[301];
assign xnor7[302] = 1'b1 ^~ inbuffer_data[302];
assign xnor7[303] = 1'b0 ^~ inbuffer_data[303];
assign xnor7[304] = 1'b0 ^~ inbuffer_data[304];
assign xnor7[305] = 1'b0 ^~ inbuffer_data[305];
assign xnor7[306] = 1'b1 ^~ inbuffer_data[306];
assign xnor7[307] = 1'b0 ^~ inbuffer_data[307];
assign xnor7[308] = 1'b0 ^~ inbuffer_data[308];
assign xnor7[309] = 1'b1 ^~ inbuffer_data[309];
assign xnor7[310] = 1'b1 ^~ inbuffer_data[310];
assign xnor7[311] = 1'b1 ^~ inbuffer_data[311];
assign xnor7[312] = 1'b1 ^~ inbuffer_data[312];
assign xnor7[313] = 1'b1 ^~ inbuffer_data[313];
assign xnor7[314] = 1'b1 ^~ inbuffer_data[314];
assign xnor7[315] = 1'b1 ^~ inbuffer_data[315];
assign xnor7[316] = 1'b1 ^~ inbuffer_data[316];
assign xnor7[317] = 1'b1 ^~ inbuffer_data[317];
assign xnor7[318] = 1'b1 ^~ inbuffer_data[318];
assign xnor7[319] = 1'b0 ^~ inbuffer_data[319];
assign xnor7[320] = 1'b0 ^~ inbuffer_data[320];
assign xnor7[321] = 1'b0 ^~ inbuffer_data[321];
assign xnor7[322] = 1'b1 ^~ inbuffer_data[322];
assign xnor7[323] = 1'b1 ^~ inbuffer_data[323];
assign xnor7[324] = 1'b1 ^~ inbuffer_data[324];
assign xnor7[325] = 1'b1 ^~ inbuffer_data[325];
assign xnor7[326] = 1'b1 ^~ inbuffer_data[326];
assign xnor7[327] = 1'b1 ^~ inbuffer_data[327];
assign xnor7[328] = 1'b1 ^~ inbuffer_data[328];
assign xnor7[329] = 1'b1 ^~ inbuffer_data[329];
assign xnor7[330] = 1'b1 ^~ inbuffer_data[330];
assign xnor7[331] = 1'b0 ^~ inbuffer_data[331];
assign xnor7[332] = 1'b0 ^~ inbuffer_data[332];
assign xnor7[333] = 1'b0 ^~ inbuffer_data[333];
assign xnor7[334] = 1'b0 ^~ inbuffer_data[334];
assign xnor7[335] = 1'b0 ^~ inbuffer_data[335];
assign xnor7[336] = 1'b0 ^~ inbuffer_data[336];
assign xnor7[337] = 1'b0 ^~ inbuffer_data[337];
assign xnor7[338] = 1'b1 ^~ inbuffer_data[338];
assign xnor7[339] = 1'b1 ^~ inbuffer_data[339];
assign xnor7[340] = 1'b1 ^~ inbuffer_data[340];
assign xnor7[341] = 1'b1 ^~ inbuffer_data[341];
assign xnor7[342] = 1'b1 ^~ inbuffer_data[342];
assign xnor7[343] = 1'b1 ^~ inbuffer_data[343];
assign xnor7[344] = 1'b1 ^~ inbuffer_data[344];
assign xnor7[345] = 1'b1 ^~ inbuffer_data[345];
assign xnor7[346] = 1'b0 ^~ inbuffer_data[346];
assign xnor7[347] = 1'b0 ^~ inbuffer_data[347];
assign xnor7[348] = 1'b0 ^~ inbuffer_data[348];
assign xnor7[349] = 1'b0 ^~ inbuffer_data[349];
assign xnor7[350] = 1'b0 ^~ inbuffer_data[350];
assign xnor7[351] = 1'b1 ^~ inbuffer_data[351];
assign xnor7[352] = 1'b1 ^~ inbuffer_data[352];
assign xnor7[353] = 1'b1 ^~ inbuffer_data[353];
assign xnor7[354] = 1'b1 ^~ inbuffer_data[354];
assign xnor7[355] = 1'b0 ^~ inbuffer_data[355];
assign xnor7[356] = 1'b0 ^~ inbuffer_data[356];
assign xnor7[357] = 1'b0 ^~ inbuffer_data[357];
assign xnor7[358] = 1'b1 ^~ inbuffer_data[358];
assign xnor7[359] = 1'b0 ^~ inbuffer_data[359];
assign xnor7[360] = 1'b0 ^~ inbuffer_data[360];
assign xnor7[361] = 1'b0 ^~ inbuffer_data[361];
assign xnor7[362] = 1'b0 ^~ inbuffer_data[362];
assign xnor7[363] = 1'b1 ^~ inbuffer_data[363];
assign xnor7[364] = 1'b0 ^~ inbuffer_data[364];
assign xnor7[365] = 1'b1 ^~ inbuffer_data[365];
assign xnor7[366] = 1'b1 ^~ inbuffer_data[366];
assign xnor7[367] = 1'b1 ^~ inbuffer_data[367];
assign xnor7[368] = 1'b1 ^~ inbuffer_data[368];
assign xnor7[369] = 1'b1 ^~ inbuffer_data[369];
assign xnor7[370] = 1'b1 ^~ inbuffer_data[370];
assign xnor7[371] = 1'b1 ^~ inbuffer_data[371];
assign xnor7[372] = 1'b0 ^~ inbuffer_data[372];
assign xnor7[373] = 1'b0 ^~ inbuffer_data[373];
assign xnor7[374] = 1'b0 ^~ inbuffer_data[374];
assign xnor7[375] = 1'b0 ^~ inbuffer_data[375];
assign xnor7[376] = 1'b0 ^~ inbuffer_data[376];
assign xnor7[377] = 1'b0 ^~ inbuffer_data[377];
assign xnor7[378] = 1'b0 ^~ inbuffer_data[378];
assign xnor7[379] = 1'b1 ^~ inbuffer_data[379];
assign xnor7[380] = 1'b1 ^~ inbuffer_data[380];
assign xnor7[381] = 1'b1 ^~ inbuffer_data[381];
assign xnor7[382] = 1'b0 ^~ inbuffer_data[382];
assign xnor7[383] = 1'b0 ^~ inbuffer_data[383];
assign xnor7[384] = 1'b1 ^~ inbuffer_data[384];
assign xnor7[385] = 1'b0 ^~ inbuffer_data[385];
assign xnor7[386] = 1'b0 ^~ inbuffer_data[386];
assign xnor7[387] = 1'b0 ^~ inbuffer_data[387];
assign xnor7[388] = 1'b1 ^~ inbuffer_data[388];
assign xnor7[389] = 1'b1 ^~ inbuffer_data[389];
assign xnor7[390] = 1'b0 ^~ inbuffer_data[390];
assign xnor7[391] = 1'b0 ^~ inbuffer_data[391];
assign xnor7[392] = 1'b0 ^~ inbuffer_data[392];
assign xnor7[393] = 1'b1 ^~ inbuffer_data[393];
assign xnor7[394] = 1'b0 ^~ inbuffer_data[394];
assign xnor7[395] = 1'b0 ^~ inbuffer_data[395];
assign xnor7[396] = 1'b0 ^~ inbuffer_data[396];
assign xnor7[397] = 1'b1 ^~ inbuffer_data[397];
assign xnor7[398] = 1'b0 ^~ inbuffer_data[398];
assign xnor7[399] = 1'b1 ^~ inbuffer_data[399];
assign xnor7[400] = 1'b0 ^~ inbuffer_data[400];
assign xnor7[401] = 1'b0 ^~ inbuffer_data[401];
assign xnor7[402] = 1'b0 ^~ inbuffer_data[402];
assign xnor7[403] = 1'b0 ^~ inbuffer_data[403];
assign xnor7[404] = 1'b0 ^~ inbuffer_data[404];
assign xnor7[405] = 1'b0 ^~ inbuffer_data[405];
assign xnor7[406] = 1'b0 ^~ inbuffer_data[406];
assign xnor7[407] = 1'b1 ^~ inbuffer_data[407];
assign xnor7[408] = 1'b1 ^~ inbuffer_data[408];
assign xnor7[409] = 1'b1 ^~ inbuffer_data[409];
assign xnor7[410] = 1'b1 ^~ inbuffer_data[410];
assign xnor7[411] = 1'b1 ^~ inbuffer_data[411];
assign xnor7[412] = 1'b1 ^~ inbuffer_data[412];
assign xnor7[413] = 1'b1 ^~ inbuffer_data[413];
assign xnor7[414] = 1'b1 ^~ inbuffer_data[414];
assign xnor7[415] = 1'b1 ^~ inbuffer_data[415];
assign xnor7[416] = 1'b0 ^~ inbuffer_data[416];
assign xnor7[417] = 1'b0 ^~ inbuffer_data[417];
assign xnor7[418] = 1'b0 ^~ inbuffer_data[418];
assign xnor7[419] = 1'b0 ^~ inbuffer_data[419];
assign xnor7[420] = 1'b1 ^~ inbuffer_data[420];
assign xnor7[421] = 1'b1 ^~ inbuffer_data[421];
assign xnor7[422] = 1'b0 ^~ inbuffer_data[422];
assign xnor7[423] = 1'b1 ^~ inbuffer_data[423];
assign xnor7[424] = 1'b0 ^~ inbuffer_data[424];
assign xnor7[425] = 1'b1 ^~ inbuffer_data[425];
assign xnor7[426] = 1'b1 ^~ inbuffer_data[426];
assign xnor7[427] = 1'b0 ^~ inbuffer_data[427];
assign xnor7[428] = 1'b0 ^~ inbuffer_data[428];
assign xnor7[429] = 1'b0 ^~ inbuffer_data[429];
assign xnor7[430] = 1'b0 ^~ inbuffer_data[430];
assign xnor7[431] = 1'b0 ^~ inbuffer_data[431];
assign xnor7[432] = 1'b0 ^~ inbuffer_data[432];
assign xnor7[433] = 1'b0 ^~ inbuffer_data[433];
assign xnor7[434] = 1'b0 ^~ inbuffer_data[434];
assign xnor7[435] = 1'b0 ^~ inbuffer_data[435];
assign xnor7[436] = 1'b0 ^~ inbuffer_data[436];
assign xnor7[437] = 1'b1 ^~ inbuffer_data[437];
assign xnor7[438] = 1'b1 ^~ inbuffer_data[438];
assign xnor7[439] = 1'b1 ^~ inbuffer_data[439];
assign xnor7[440] = 1'b1 ^~ inbuffer_data[440];
assign xnor7[441] = 1'b1 ^~ inbuffer_data[441];
assign xnor7[442] = 1'b1 ^~ inbuffer_data[442];
assign xnor7[443] = 1'b1 ^~ inbuffer_data[443];
assign xnor7[444] = 1'b1 ^~ inbuffer_data[444];
assign xnor7[445] = 1'b1 ^~ inbuffer_data[445];
assign xnor7[446] = 1'b0 ^~ inbuffer_data[446];
assign xnor7[447] = 1'b0 ^~ inbuffer_data[447];
assign xnor7[448] = 1'b1 ^~ inbuffer_data[448];
assign xnor7[449] = 1'b1 ^~ inbuffer_data[449];
assign xnor7[450] = 1'b1 ^~ inbuffer_data[450];
assign xnor7[451] = 1'b0 ^~ inbuffer_data[451];
assign xnor7[452] = 1'b1 ^~ inbuffer_data[452];
assign xnor7[453] = 1'b0 ^~ inbuffer_data[453];
assign xnor7[454] = 1'b1 ^~ inbuffer_data[454];
assign xnor7[455] = 1'b1 ^~ inbuffer_data[455];
assign xnor7[456] = 1'b1 ^~ inbuffer_data[456];
assign xnor7[457] = 1'b0 ^~ inbuffer_data[457];
assign xnor7[458] = 1'b0 ^~ inbuffer_data[458];
assign xnor7[459] = 1'b0 ^~ inbuffer_data[459];
assign xnor7[460] = 1'b0 ^~ inbuffer_data[460];
assign xnor7[461] = 1'b0 ^~ inbuffer_data[461];
assign xnor7[462] = 1'b0 ^~ inbuffer_data[462];
assign xnor7[463] = 1'b1 ^~ inbuffer_data[463];
assign xnor7[464] = 1'b1 ^~ inbuffer_data[464];
assign xnor7[465] = 1'b1 ^~ inbuffer_data[465];
assign xnor7[466] = 1'b1 ^~ inbuffer_data[466];
assign xnor7[467] = 1'b1 ^~ inbuffer_data[467];
assign xnor7[468] = 1'b1 ^~ inbuffer_data[468];
assign xnor7[469] = 1'b1 ^~ inbuffer_data[469];
assign xnor7[470] = 1'b0 ^~ inbuffer_data[470];
assign xnor7[471] = 1'b0 ^~ inbuffer_data[471];
assign xnor7[472] = 1'b0 ^~ inbuffer_data[472];
assign xnor7[473] = 1'b0 ^~ inbuffer_data[473];
assign xnor7[474] = 1'b0 ^~ inbuffer_data[474];
assign xnor7[475] = 1'b1 ^~ inbuffer_data[475];
assign xnor7[476] = 1'b0 ^~ inbuffer_data[476];
assign xnor7[477] = 1'b1 ^~ inbuffer_data[477];
assign xnor7[478] = 1'b1 ^~ inbuffer_data[478];
assign xnor7[479] = 1'b0 ^~ inbuffer_data[479];
assign xnor7[480] = 1'b1 ^~ inbuffer_data[480];
assign xnor7[481] = 1'b0 ^~ inbuffer_data[481];
assign xnor7[482] = 1'b0 ^~ inbuffer_data[482];
assign xnor7[483] = 1'b0 ^~ inbuffer_data[483];
assign xnor7[484] = 1'b0 ^~ inbuffer_data[484];
assign xnor7[485] = 1'b0 ^~ inbuffer_data[485];
assign xnor7[486] = 1'b0 ^~ inbuffer_data[486];
assign xnor7[487] = 1'b0 ^~ inbuffer_data[487];
assign xnor7[488] = 1'b1 ^~ inbuffer_data[488];
assign xnor7[489] = 1'b1 ^~ inbuffer_data[489];
assign xnor7[490] = 1'b1 ^~ inbuffer_data[490];
assign xnor7[491] = 1'b1 ^~ inbuffer_data[491];
assign xnor7[492] = 1'b1 ^~ inbuffer_data[492];
assign xnor7[493] = 1'b1 ^~ inbuffer_data[493];
assign xnor7[494] = 1'b1 ^~ inbuffer_data[494];
assign xnor7[495] = 1'b0 ^~ inbuffer_data[495];
assign xnor7[496] = 1'b1 ^~ inbuffer_data[496];
assign xnor7[497] = 1'b1 ^~ inbuffer_data[497];
assign xnor7[498] = 1'b0 ^~ inbuffer_data[498];
assign xnor7[499] = 1'b0 ^~ inbuffer_data[499];
assign xnor7[500] = 1'b1 ^~ inbuffer_data[500];
assign xnor7[501] = 1'b0 ^~ inbuffer_data[501];
assign xnor7[502] = 1'b1 ^~ inbuffer_data[502];
assign xnor7[503] = 1'b1 ^~ inbuffer_data[503];
assign xnor7[504] = 1'b0 ^~ inbuffer_data[504];
assign xnor7[505] = 1'b1 ^~ inbuffer_data[505];
assign xnor7[506] = 1'b0 ^~ inbuffer_data[506];
assign xnor7[507] = 1'b0 ^~ inbuffer_data[507];
assign xnor7[508] = 1'b1 ^~ inbuffer_data[508];
assign xnor7[509] = 1'b0 ^~ inbuffer_data[509];
assign xnor7[510] = 1'b0 ^~ inbuffer_data[510];
assign xnor7[511] = 1'b0 ^~ inbuffer_data[511];
assign xnor7[512] = 1'b0 ^~ inbuffer_data[512];
assign xnor7[513] = 1'b0 ^~ inbuffer_data[513];
assign xnor7[514] = 1'b0 ^~ inbuffer_data[514];
assign xnor7[515] = 1'b0 ^~ inbuffer_data[515];
assign xnor7[516] = 1'b0 ^~ inbuffer_data[516];
assign xnor7[517] = 1'b1 ^~ inbuffer_data[517];
assign xnor7[518] = 1'b1 ^~ inbuffer_data[518];
assign xnor7[519] = 1'b1 ^~ inbuffer_data[519];
assign xnor7[520] = 1'b1 ^~ inbuffer_data[520];
assign xnor7[521] = 1'b0 ^~ inbuffer_data[521];
assign xnor7[522] = 1'b0 ^~ inbuffer_data[522];
assign xnor7[523] = 1'b1 ^~ inbuffer_data[523];
assign xnor7[524] = 1'b0 ^~ inbuffer_data[524];
assign xnor7[525] = 1'b0 ^~ inbuffer_data[525];
assign xnor7[526] = 1'b0 ^~ inbuffer_data[526];
assign xnor7[527] = 1'b0 ^~ inbuffer_data[527];
assign xnor7[528] = 1'b0 ^~ inbuffer_data[528];
assign xnor7[529] = 1'b0 ^~ inbuffer_data[529];
assign xnor7[530] = 1'b0 ^~ inbuffer_data[530];
assign xnor7[531] = 1'b1 ^~ inbuffer_data[531];
assign xnor7[532] = 1'b1 ^~ inbuffer_data[532];
assign xnor7[533] = 1'b1 ^~ inbuffer_data[533];
assign xnor7[534] = 1'b1 ^~ inbuffer_data[534];
assign xnor7[535] = 1'b1 ^~ inbuffer_data[535];
assign xnor7[536] = 1'b1 ^~ inbuffer_data[536];
assign xnor7[537] = 1'b0 ^~ inbuffer_data[537];
assign xnor7[538] = 1'b0 ^~ inbuffer_data[538];
assign xnor7[539] = 1'b0 ^~ inbuffer_data[539];
assign xnor7[540] = 1'b0 ^~ inbuffer_data[540];
assign xnor7[541] = 1'b0 ^~ inbuffer_data[541];
assign xnor7[542] = 1'b0 ^~ inbuffer_data[542];
assign xnor7[543] = 1'b0 ^~ inbuffer_data[543];
assign xnor7[544] = 1'b1 ^~ inbuffer_data[544];
assign xnor7[545] = 1'b0 ^~ inbuffer_data[545];
assign xnor7[546] = 1'b1 ^~ inbuffer_data[546];
assign xnor7[547] = 1'b0 ^~ inbuffer_data[547];
assign xnor7[548] = 1'b0 ^~ inbuffer_data[548];
assign xnor7[549] = 1'b0 ^~ inbuffer_data[549];
assign xnor7[550] = 1'b0 ^~ inbuffer_data[550];
assign xnor7[551] = 1'b0 ^~ inbuffer_data[551];
assign xnor7[552] = 1'b0 ^~ inbuffer_data[552];
assign xnor7[553] = 1'b0 ^~ inbuffer_data[553];
assign xnor7[554] = 1'b0 ^~ inbuffer_data[554];
assign xnor7[555] = 1'b0 ^~ inbuffer_data[555];
assign xnor7[556] = 1'b0 ^~ inbuffer_data[556];
assign xnor7[557] = 1'b0 ^~ inbuffer_data[557];
assign xnor7[558] = 1'b0 ^~ inbuffer_data[558];
assign xnor7[559] = 1'b1 ^~ inbuffer_data[559];
assign xnor7[560] = 1'b1 ^~ inbuffer_data[560];
assign xnor7[561] = 1'b0 ^~ inbuffer_data[561];
assign xnor7[562] = 1'b0 ^~ inbuffer_data[562];
assign xnor7[563] = 1'b0 ^~ inbuffer_data[563];
assign xnor7[564] = 1'b0 ^~ inbuffer_data[564];
assign xnor7[565] = 1'b0 ^~ inbuffer_data[565];
assign xnor7[566] = 1'b0 ^~ inbuffer_data[566];
assign xnor7[567] = 1'b0 ^~ inbuffer_data[567];
assign xnor7[568] = 1'b0 ^~ inbuffer_data[568];
assign xnor7[569] = 1'b0 ^~ inbuffer_data[569];
assign xnor7[570] = 1'b0 ^~ inbuffer_data[570];
assign xnor7[571] = 1'b1 ^~ inbuffer_data[571];
assign xnor7[572] = 1'b1 ^~ inbuffer_data[572];
assign xnor7[573] = 1'b1 ^~ inbuffer_data[573];
assign xnor7[574] = 1'b1 ^~ inbuffer_data[574];
assign xnor7[575] = 1'b0 ^~ inbuffer_data[575];
assign xnor7[576] = 1'b0 ^~ inbuffer_data[576];
assign xnor7[577] = 1'b0 ^~ inbuffer_data[577];
assign xnor7[578] = 1'b0 ^~ inbuffer_data[578];
assign xnor7[579] = 1'b0 ^~ inbuffer_data[579];
assign xnor7[580] = 1'b0 ^~ inbuffer_data[580];
assign xnor7[581] = 1'b0 ^~ inbuffer_data[581];
assign xnor7[582] = 1'b0 ^~ inbuffer_data[582];
assign xnor7[583] = 1'b0 ^~ inbuffer_data[583];
assign xnor7[584] = 1'b0 ^~ inbuffer_data[584];
assign xnor7[585] = 1'b0 ^~ inbuffer_data[585];
assign xnor7[586] = 1'b1 ^~ inbuffer_data[586];
assign xnor7[587] = 1'b1 ^~ inbuffer_data[587];
assign xnor7[588] = 1'b0 ^~ inbuffer_data[588];
assign xnor7[589] = 1'b1 ^~ inbuffer_data[589];
assign xnor7[590] = 1'b0 ^~ inbuffer_data[590];
assign xnor7[591] = 1'b0 ^~ inbuffer_data[591];
assign xnor7[592] = 1'b0 ^~ inbuffer_data[592];
assign xnor7[593] = 1'b0 ^~ inbuffer_data[593];
assign xnor7[594] = 1'b0 ^~ inbuffer_data[594];
assign xnor7[595] = 1'b0 ^~ inbuffer_data[595];
assign xnor7[596] = 1'b0 ^~ inbuffer_data[596];
assign xnor7[597] = 1'b0 ^~ inbuffer_data[597];
assign xnor7[598] = 1'b1 ^~ inbuffer_data[598];
assign xnor7[599] = 1'b0 ^~ inbuffer_data[599];
assign xnor7[600] = 1'b0 ^~ inbuffer_data[600];
assign xnor7[601] = 1'b0 ^~ inbuffer_data[601];
assign xnor7[602] = 1'b0 ^~ inbuffer_data[602];
assign xnor7[603] = 1'b0 ^~ inbuffer_data[603];
assign xnor7[604] = 1'b0 ^~ inbuffer_data[604];
assign xnor7[605] = 1'b0 ^~ inbuffer_data[605];
assign xnor7[606] = 1'b0 ^~ inbuffer_data[606];
assign xnor7[607] = 1'b0 ^~ inbuffer_data[607];
assign xnor7[608] = 1'b0 ^~ inbuffer_data[608];
assign xnor7[609] = 1'b0 ^~ inbuffer_data[609];
assign xnor7[610] = 1'b0 ^~ inbuffer_data[610];
assign xnor7[611] = 1'b0 ^~ inbuffer_data[611];
assign xnor7[612] = 1'b1 ^~ inbuffer_data[612];
assign xnor7[613] = 1'b1 ^~ inbuffer_data[613];
assign xnor7[614] = 1'b0 ^~ inbuffer_data[614];
assign xnor7[615] = 1'b0 ^~ inbuffer_data[615];
assign xnor7[616] = 1'b1 ^~ inbuffer_data[616];
assign xnor7[617] = 1'b1 ^~ inbuffer_data[617];
assign xnor7[618] = 1'b1 ^~ inbuffer_data[618];
assign xnor7[619] = 1'b1 ^~ inbuffer_data[619];
assign xnor7[620] = 1'b0 ^~ inbuffer_data[620];
assign xnor7[621] = 1'b0 ^~ inbuffer_data[621];
assign xnor7[622] = 1'b0 ^~ inbuffer_data[622];
assign xnor7[623] = 1'b1 ^~ inbuffer_data[623];
assign xnor7[624] = 1'b1 ^~ inbuffer_data[624];
assign xnor7[625] = 1'b1 ^~ inbuffer_data[625];
assign xnor7[626] = 1'b0 ^~ inbuffer_data[626];
assign xnor7[627] = 1'b0 ^~ inbuffer_data[627];
assign xnor7[628] = 1'b0 ^~ inbuffer_data[628];
assign xnor7[629] = 1'b0 ^~ inbuffer_data[629];
assign xnor7[630] = 1'b0 ^~ inbuffer_data[630];
assign xnor7[631] = 1'b0 ^~ inbuffer_data[631];
assign xnor7[632] = 1'b0 ^~ inbuffer_data[632];
assign xnor7[633] = 1'b0 ^~ inbuffer_data[633];
assign xnor7[634] = 1'b0 ^~ inbuffer_data[634];
assign xnor7[635] = 1'b0 ^~ inbuffer_data[635];
assign xnor7[636] = 1'b0 ^~ inbuffer_data[636];
assign xnor7[637] = 1'b0 ^~ inbuffer_data[637];
assign xnor7[638] = 1'b0 ^~ inbuffer_data[638];
assign xnor7[639] = 1'b0 ^~ inbuffer_data[639];
assign xnor7[640] = 1'b0 ^~ inbuffer_data[640];
assign xnor7[641] = 1'b1 ^~ inbuffer_data[641];
assign xnor7[642] = 1'b0 ^~ inbuffer_data[642];
assign xnor7[643] = 1'b1 ^~ inbuffer_data[643];
assign xnor7[644] = 1'b1 ^~ inbuffer_data[644];
assign xnor7[645] = 1'b0 ^~ inbuffer_data[645];
assign xnor7[646] = 1'b1 ^~ inbuffer_data[646];
assign xnor7[647] = 1'b0 ^~ inbuffer_data[647];
assign xnor7[648] = 1'b0 ^~ inbuffer_data[648];
assign xnor7[649] = 1'b1 ^~ inbuffer_data[649];
assign xnor7[650] = 1'b1 ^~ inbuffer_data[650];
assign xnor7[651] = 1'b1 ^~ inbuffer_data[651];
assign xnor7[652] = 1'b0 ^~ inbuffer_data[652];
assign xnor7[653] = 1'b0 ^~ inbuffer_data[653];
assign xnor7[654] = 1'b0 ^~ inbuffer_data[654];
assign xnor7[655] = 1'b1 ^~ inbuffer_data[655];
assign xnor7[656] = 1'b0 ^~ inbuffer_data[656];
assign xnor7[657] = 1'b0 ^~ inbuffer_data[657];
assign xnor7[658] = 1'b0 ^~ inbuffer_data[658];
assign xnor7[659] = 1'b1 ^~ inbuffer_data[659];
assign xnor7[660] = 1'b1 ^~ inbuffer_data[660];
assign xnor7[661] = 1'b1 ^~ inbuffer_data[661];
assign xnor7[662] = 1'b0 ^~ inbuffer_data[662];
assign xnor7[663] = 1'b0 ^~ inbuffer_data[663];
assign xnor7[664] = 1'b0 ^~ inbuffer_data[664];
assign xnor7[665] = 1'b0 ^~ inbuffer_data[665];
assign xnor7[666] = 1'b0 ^~ inbuffer_data[666];
assign xnor7[667] = 1'b0 ^~ inbuffer_data[667];
assign xnor7[668] = 1'b1 ^~ inbuffer_data[668];
assign xnor7[669] = 1'b0 ^~ inbuffer_data[669];
assign xnor7[670] = 1'b1 ^~ inbuffer_data[670];
assign xnor7[671] = 1'b1 ^~ inbuffer_data[671];
assign xnor7[672] = 1'b1 ^~ inbuffer_data[672];
assign xnor7[673] = 1'b1 ^~ inbuffer_data[673];
assign xnor7[674] = 1'b0 ^~ inbuffer_data[674];
assign xnor7[675] = 1'b1 ^~ inbuffer_data[675];
assign xnor7[676] = 1'b0 ^~ inbuffer_data[676];
assign xnor7[677] = 1'b1 ^~ inbuffer_data[677];
assign xnor7[678] = 1'b1 ^~ inbuffer_data[678];
assign xnor7[679] = 1'b1 ^~ inbuffer_data[679];
assign xnor7[680] = 1'b1 ^~ inbuffer_data[680];
assign xnor7[681] = 1'b0 ^~ inbuffer_data[681];
assign xnor7[682] = 1'b1 ^~ inbuffer_data[682];
assign xnor7[683] = 1'b1 ^~ inbuffer_data[683];
assign xnor7[684] = 1'b1 ^~ inbuffer_data[684];
assign xnor7[685] = 1'b1 ^~ inbuffer_data[685];
assign xnor7[686] = 1'b1 ^~ inbuffer_data[686];
assign xnor7[687] = 1'b0 ^~ inbuffer_data[687];
assign xnor7[688] = 1'b1 ^~ inbuffer_data[688];
assign xnor7[689] = 1'b0 ^~ inbuffer_data[689];
assign xnor7[690] = 1'b0 ^~ inbuffer_data[690];
assign xnor7[691] = 1'b0 ^~ inbuffer_data[691];
assign xnor7[692] = 1'b0 ^~ inbuffer_data[692];
assign xnor7[693] = 1'b0 ^~ inbuffer_data[693];
assign xnor7[694] = 1'b0 ^~ inbuffer_data[694];
assign xnor7[695] = 1'b0 ^~ inbuffer_data[695];
assign xnor7[696] = 1'b1 ^~ inbuffer_data[696];
assign xnor7[697] = 1'b1 ^~ inbuffer_data[697];
assign xnor7[698] = 1'b1 ^~ inbuffer_data[698];
assign xnor7[699] = 1'b0 ^~ inbuffer_data[699];
assign xnor7[700] = 1'b0 ^~ inbuffer_data[700];
assign xnor7[701] = 1'b0 ^~ inbuffer_data[701];
assign xnor7[702] = 1'b1 ^~ inbuffer_data[702];
assign xnor7[703] = 1'b0 ^~ inbuffer_data[703];
assign xnor7[704] = 1'b1 ^~ inbuffer_data[704];
assign xnor7[705] = 1'b0 ^~ inbuffer_data[705];
assign xnor7[706] = 1'b0 ^~ inbuffer_data[706];
assign xnor7[707] = 1'b1 ^~ inbuffer_data[707];
assign xnor7[708] = 1'b1 ^~ inbuffer_data[708];
assign xnor7[709] = 1'b1 ^~ inbuffer_data[709];
assign xnor7[710] = 1'b1 ^~ inbuffer_data[710];
assign xnor7[711] = 1'b1 ^~ inbuffer_data[711];
assign xnor7[712] = 1'b1 ^~ inbuffer_data[712];
assign xnor7[713] = 1'b1 ^~ inbuffer_data[713];
assign xnor7[714] = 1'b1 ^~ inbuffer_data[714];
assign xnor7[715] = 1'b1 ^~ inbuffer_data[715];
assign xnor7[716] = 1'b1 ^~ inbuffer_data[716];
assign xnor7[717] = 1'b1 ^~ inbuffer_data[717];
assign xnor7[718] = 1'b1 ^~ inbuffer_data[718];
assign xnor7[719] = 1'b1 ^~ inbuffer_data[719];
assign xnor7[720] = 1'b1 ^~ inbuffer_data[720];
assign xnor7[721] = 1'b0 ^~ inbuffer_data[721];
assign xnor7[722] = 1'b1 ^~ inbuffer_data[722];
assign xnor7[723] = 1'b0 ^~ inbuffer_data[723];
assign xnor7[724] = 1'b1 ^~ inbuffer_data[724];
assign xnor7[725] = 1'b0 ^~ inbuffer_data[725];
assign xnor7[726] = 1'b0 ^~ inbuffer_data[726];
assign xnor7[727] = 1'b1 ^~ inbuffer_data[727];
assign xnor7[728] = 1'b0 ^~ inbuffer_data[728];
assign xnor7[729] = 1'b0 ^~ inbuffer_data[729];
assign xnor7[730] = 1'b1 ^~ inbuffer_data[730];
assign xnor7[731] = 1'b1 ^~ inbuffer_data[731];
assign xnor7[732] = 1'b1 ^~ inbuffer_data[732];
assign xnor7[733] = 1'b1 ^~ inbuffer_data[733];
assign xnor7[734] = 1'b0 ^~ inbuffer_data[734];
assign xnor7[735] = 1'b1 ^~ inbuffer_data[735];
assign xnor7[736] = 1'b1 ^~ inbuffer_data[736];
assign xnor7[737] = 1'b1 ^~ inbuffer_data[737];
assign xnor7[738] = 1'b1 ^~ inbuffer_data[738];
assign xnor7[739] = 1'b0 ^~ inbuffer_data[739];
assign xnor7[740] = 1'b1 ^~ inbuffer_data[740];
assign xnor7[741] = 1'b1 ^~ inbuffer_data[741];
assign xnor7[742] = 1'b1 ^~ inbuffer_data[742];
assign xnor7[743] = 1'b1 ^~ inbuffer_data[743];
assign xnor7[744] = 1'b1 ^~ inbuffer_data[744];
assign xnor7[745] = 1'b1 ^~ inbuffer_data[745];
assign xnor7[746] = 1'b1 ^~ inbuffer_data[746];
assign xnor7[747] = 1'b1 ^~ inbuffer_data[747];
assign xnor7[748] = 1'b0 ^~ inbuffer_data[748];
assign xnor7[749] = 1'b1 ^~ inbuffer_data[749];
assign xnor7[750] = 1'b0 ^~ inbuffer_data[750];
assign xnor7[751] = 1'b0 ^~ inbuffer_data[751];
assign xnor7[752] = 1'b0 ^~ inbuffer_data[752];
assign xnor7[753] = 1'b1 ^~ inbuffer_data[753];
assign xnor7[754] = 1'b1 ^~ inbuffer_data[754];
assign xnor7[755] = 1'b0 ^~ inbuffer_data[755];
assign xnor7[756] = 1'b1 ^~ inbuffer_data[756];
assign xnor7[757] = 1'b0 ^~ inbuffer_data[757];
assign xnor7[758] = 1'b1 ^~ inbuffer_data[758];
assign xnor7[759] = 1'b0 ^~ inbuffer_data[759];
assign xnor7[760] = 1'b0 ^~ inbuffer_data[760];
assign xnor7[761] = 1'b1 ^~ inbuffer_data[761];
assign xnor7[762] = 1'b1 ^~ inbuffer_data[762];
assign xnor7[763] = 1'b0 ^~ inbuffer_data[763];
assign xnor7[764] = 1'b0 ^~ inbuffer_data[764];
assign xnor7[765] = 1'b1 ^~ inbuffer_data[765];
assign xnor7[766] = 1'b0 ^~ inbuffer_data[766];
assign xnor7[767] = 1'b0 ^~ inbuffer_data[767];
assign xnor7[768] = 1'b0 ^~ inbuffer_data[768];
assign xnor7[769] = 1'b0 ^~ inbuffer_data[769];
assign xnor7[770] = 1'b1 ^~ inbuffer_data[770];
assign xnor7[771] = 1'b1 ^~ inbuffer_data[771];
assign xnor7[772] = 1'b1 ^~ inbuffer_data[772];
assign xnor7[773] = 1'b0 ^~ inbuffer_data[773];
assign xnor7[774] = 1'b0 ^~ inbuffer_data[774];
assign xnor7[775] = 1'b1 ^~ inbuffer_data[775];
assign xnor7[776] = 1'b1 ^~ inbuffer_data[776];
assign xnor7[777] = 1'b0 ^~ inbuffer_data[777];
assign xnor7[778] = 1'b1 ^~ inbuffer_data[778];
assign xnor7[779] = 1'b0 ^~ inbuffer_data[779];
assign xnor7[780] = 1'b1 ^~ inbuffer_data[780];
assign xnor7[781] = 1'b0 ^~ inbuffer_data[781];
assign xnor7[782] = 1'b0 ^~ inbuffer_data[782];
assign xnor7[783] = 1'b1 ^~ inbuffer_data[783];
assign xnor8[0] = 1'b1 ^~ inbuffer_data[0];
assign xnor8[1] = 1'b1 ^~ inbuffer_data[1];
assign xnor8[2] = 1'b1 ^~ inbuffer_data[2];
assign xnor8[3] = 1'b1 ^~ inbuffer_data[3];
assign xnor8[4] = 1'b1 ^~ inbuffer_data[4];
assign xnor8[5] = 1'b0 ^~ inbuffer_data[5];
assign xnor8[6] = 1'b0 ^~ inbuffer_data[6];
assign xnor8[7] = 1'b0 ^~ inbuffer_data[7];
assign xnor8[8] = 1'b1 ^~ inbuffer_data[8];
assign xnor8[9] = 1'b0 ^~ inbuffer_data[9];
assign xnor8[10] = 1'b1 ^~ inbuffer_data[10];
assign xnor8[11] = 1'b0 ^~ inbuffer_data[11];
assign xnor8[12] = 1'b0 ^~ inbuffer_data[12];
assign xnor8[13] = 1'b0 ^~ inbuffer_data[13];
assign xnor8[14] = 1'b1 ^~ inbuffer_data[14];
assign xnor8[15] = 1'b1 ^~ inbuffer_data[15];
assign xnor8[16] = 1'b0 ^~ inbuffer_data[16];
assign xnor8[17] = 1'b1 ^~ inbuffer_data[17];
assign xnor8[18] = 1'b0 ^~ inbuffer_data[18];
assign xnor8[19] = 1'b0 ^~ inbuffer_data[19];
assign xnor8[20] = 1'b0 ^~ inbuffer_data[20];
assign xnor8[21] = 1'b1 ^~ inbuffer_data[21];
assign xnor8[22] = 1'b0 ^~ inbuffer_data[22];
assign xnor8[23] = 1'b1 ^~ inbuffer_data[23];
assign xnor8[24] = 1'b1 ^~ inbuffer_data[24];
assign xnor8[25] = 1'b1 ^~ inbuffer_data[25];
assign xnor8[26] = 1'b1 ^~ inbuffer_data[26];
assign xnor8[27] = 1'b0 ^~ inbuffer_data[27];
assign xnor8[28] = 1'b1 ^~ inbuffer_data[28];
assign xnor8[29] = 1'b1 ^~ inbuffer_data[29];
assign xnor8[30] = 1'b1 ^~ inbuffer_data[30];
assign xnor8[31] = 1'b0 ^~ inbuffer_data[31];
assign xnor8[32] = 1'b0 ^~ inbuffer_data[32];
assign xnor8[33] = 1'b1 ^~ inbuffer_data[33];
assign xnor8[34] = 1'b1 ^~ inbuffer_data[34];
assign xnor8[35] = 1'b0 ^~ inbuffer_data[35];
assign xnor8[36] = 1'b0 ^~ inbuffer_data[36];
assign xnor8[37] = 1'b0 ^~ inbuffer_data[37];
assign xnor8[38] = 1'b0 ^~ inbuffer_data[38];
assign xnor8[39] = 1'b1 ^~ inbuffer_data[39];
assign xnor8[40] = 1'b0 ^~ inbuffer_data[40];
assign xnor8[41] = 1'b1 ^~ inbuffer_data[41];
assign xnor8[42] = 1'b0 ^~ inbuffer_data[42];
assign xnor8[43] = 1'b1 ^~ inbuffer_data[43];
assign xnor8[44] = 1'b0 ^~ inbuffer_data[44];
assign xnor8[45] = 1'b0 ^~ inbuffer_data[45];
assign xnor8[46] = 1'b0 ^~ inbuffer_data[46];
assign xnor8[47] = 1'b1 ^~ inbuffer_data[47];
assign xnor8[48] = 1'b0 ^~ inbuffer_data[48];
assign xnor8[49] = 1'b1 ^~ inbuffer_data[49];
assign xnor8[50] = 1'b0 ^~ inbuffer_data[50];
assign xnor8[51] = 1'b0 ^~ inbuffer_data[51];
assign xnor8[52] = 1'b1 ^~ inbuffer_data[52];
assign xnor8[53] = 1'b0 ^~ inbuffer_data[53];
assign xnor8[54] = 1'b0 ^~ inbuffer_data[54];
assign xnor8[55] = 1'b0 ^~ inbuffer_data[55];
assign xnor8[56] = 1'b0 ^~ inbuffer_data[56];
assign xnor8[57] = 1'b1 ^~ inbuffer_data[57];
assign xnor8[58] = 1'b1 ^~ inbuffer_data[58];
assign xnor8[59] = 1'b0 ^~ inbuffer_data[59];
assign xnor8[60] = 1'b0 ^~ inbuffer_data[60];
assign xnor8[61] = 1'b0 ^~ inbuffer_data[61];
assign xnor8[62] = 1'b0 ^~ inbuffer_data[62];
assign xnor8[63] = 1'b1 ^~ inbuffer_data[63];
assign xnor8[64] = 1'b0 ^~ inbuffer_data[64];
assign xnor8[65] = 1'b1 ^~ inbuffer_data[65];
assign xnor8[66] = 1'b1 ^~ inbuffer_data[66];
assign xnor8[67] = 1'b0 ^~ inbuffer_data[67];
assign xnor8[68] = 1'b0 ^~ inbuffer_data[68];
assign xnor8[69] = 1'b0 ^~ inbuffer_data[69];
assign xnor8[70] = 1'b0 ^~ inbuffer_data[70];
assign xnor8[71] = 1'b0 ^~ inbuffer_data[71];
assign xnor8[72] = 1'b0 ^~ inbuffer_data[72];
assign xnor8[73] = 1'b0 ^~ inbuffer_data[73];
assign xnor8[74] = 1'b0 ^~ inbuffer_data[74];
assign xnor8[75] = 1'b1 ^~ inbuffer_data[75];
assign xnor8[76] = 1'b0 ^~ inbuffer_data[76];
assign xnor8[77] = 1'b0 ^~ inbuffer_data[77];
assign xnor8[78] = 1'b0 ^~ inbuffer_data[78];
assign xnor8[79] = 1'b1 ^~ inbuffer_data[79];
assign xnor8[80] = 1'b0 ^~ inbuffer_data[80];
assign xnor8[81] = 1'b1 ^~ inbuffer_data[81];
assign xnor8[82] = 1'b0 ^~ inbuffer_data[82];
assign xnor8[83] = 1'b1 ^~ inbuffer_data[83];
assign xnor8[84] = 1'b0 ^~ inbuffer_data[84];
assign xnor8[85] = 1'b0 ^~ inbuffer_data[85];
assign xnor8[86] = 1'b1 ^~ inbuffer_data[86];
assign xnor8[87] = 1'b0 ^~ inbuffer_data[87];
assign xnor8[88] = 1'b0 ^~ inbuffer_data[88];
assign xnor8[89] = 1'b1 ^~ inbuffer_data[89];
assign xnor8[90] = 1'b0 ^~ inbuffer_data[90];
assign xnor8[91] = 1'b0 ^~ inbuffer_data[91];
assign xnor8[92] = 1'b0 ^~ inbuffer_data[92];
assign xnor8[93] = 1'b0 ^~ inbuffer_data[93];
assign xnor8[94] = 1'b0 ^~ inbuffer_data[94];
assign xnor8[95] = 1'b1 ^~ inbuffer_data[95];
assign xnor8[96] = 1'b1 ^~ inbuffer_data[96];
assign xnor8[97] = 1'b0 ^~ inbuffer_data[97];
assign xnor8[98] = 1'b0 ^~ inbuffer_data[98];
assign xnor8[99] = 1'b0 ^~ inbuffer_data[99];
assign xnor8[100] = 1'b0 ^~ inbuffer_data[100];
assign xnor8[101] = 1'b0 ^~ inbuffer_data[101];
assign xnor8[102] = 1'b0 ^~ inbuffer_data[102];
assign xnor8[103] = 1'b0 ^~ inbuffer_data[103];
assign xnor8[104] = 1'b1 ^~ inbuffer_data[104];
assign xnor8[105] = 1'b1 ^~ inbuffer_data[105];
assign xnor8[106] = 1'b0 ^~ inbuffer_data[106];
assign xnor8[107] = 1'b0 ^~ inbuffer_data[107];
assign xnor8[108] = 1'b1 ^~ inbuffer_data[108];
assign xnor8[109] = 1'b0 ^~ inbuffer_data[109];
assign xnor8[110] = 1'b1 ^~ inbuffer_data[110];
assign xnor8[111] = 1'b0 ^~ inbuffer_data[111];
assign xnor8[112] = 1'b0 ^~ inbuffer_data[112];
assign xnor8[113] = 1'b1 ^~ inbuffer_data[113];
assign xnor8[114] = 1'b0 ^~ inbuffer_data[114];
assign xnor8[115] = 1'b0 ^~ inbuffer_data[115];
assign xnor8[116] = 1'b0 ^~ inbuffer_data[116];
assign xnor8[117] = 1'b0 ^~ inbuffer_data[117];
assign xnor8[118] = 1'b0 ^~ inbuffer_data[118];
assign xnor8[119] = 1'b1 ^~ inbuffer_data[119];
assign xnor8[120] = 1'b1 ^~ inbuffer_data[120];
assign xnor8[121] = 1'b0 ^~ inbuffer_data[121];
assign xnor8[122] = 1'b1 ^~ inbuffer_data[122];
assign xnor8[123] = 1'b0 ^~ inbuffer_data[123];
assign xnor8[124] = 1'b1 ^~ inbuffer_data[124];
assign xnor8[125] = 1'b1 ^~ inbuffer_data[125];
assign xnor8[126] = 1'b1 ^~ inbuffer_data[126];
assign xnor8[127] = 1'b1 ^~ inbuffer_data[127];
assign xnor8[128] = 1'b1 ^~ inbuffer_data[128];
assign xnor8[129] = 1'b1 ^~ inbuffer_data[129];
assign xnor8[130] = 1'b1 ^~ inbuffer_data[130];
assign xnor8[131] = 1'b1 ^~ inbuffer_data[131];
assign xnor8[132] = 1'b0 ^~ inbuffer_data[132];
assign xnor8[133] = 1'b1 ^~ inbuffer_data[133];
assign xnor8[134] = 1'b0 ^~ inbuffer_data[134];
assign xnor8[135] = 1'b1 ^~ inbuffer_data[135];
assign xnor8[136] = 1'b0 ^~ inbuffer_data[136];
assign xnor8[137] = 1'b0 ^~ inbuffer_data[137];
assign xnor8[138] = 1'b0 ^~ inbuffer_data[138];
assign xnor8[139] = 1'b0 ^~ inbuffer_data[139];
assign xnor8[140] = 1'b0 ^~ inbuffer_data[140];
assign xnor8[141] = 1'b0 ^~ inbuffer_data[141];
assign xnor8[142] = 1'b1 ^~ inbuffer_data[142];
assign xnor8[143] = 1'b1 ^~ inbuffer_data[143];
assign xnor8[144] = 1'b1 ^~ inbuffer_data[144];
assign xnor8[145] = 1'b0 ^~ inbuffer_data[145];
assign xnor8[146] = 1'b0 ^~ inbuffer_data[146];
assign xnor8[147] = 1'b1 ^~ inbuffer_data[147];
assign xnor8[148] = 1'b1 ^~ inbuffer_data[148];
assign xnor8[149] = 1'b1 ^~ inbuffer_data[149];
assign xnor8[150] = 1'b1 ^~ inbuffer_data[150];
assign xnor8[151] = 1'b1 ^~ inbuffer_data[151];
assign xnor8[152] = 1'b1 ^~ inbuffer_data[152];
assign xnor8[153] = 1'b1 ^~ inbuffer_data[153];
assign xnor8[154] = 1'b1 ^~ inbuffer_data[154];
assign xnor8[155] = 1'b1 ^~ inbuffer_data[155];
assign xnor8[156] = 1'b1 ^~ inbuffer_data[156];
assign xnor8[157] = 1'b1 ^~ inbuffer_data[157];
assign xnor8[158] = 1'b1 ^~ inbuffer_data[158];
assign xnor8[159] = 1'b1 ^~ inbuffer_data[159];
assign xnor8[160] = 1'b1 ^~ inbuffer_data[160];
assign xnor8[161] = 1'b1 ^~ inbuffer_data[161];
assign xnor8[162] = 1'b0 ^~ inbuffer_data[162];
assign xnor8[163] = 1'b0 ^~ inbuffer_data[163];
assign xnor8[164] = 1'b1 ^~ inbuffer_data[164];
assign xnor8[165] = 1'b0 ^~ inbuffer_data[165];
assign xnor8[166] = 1'b0 ^~ inbuffer_data[166];
assign xnor8[167] = 1'b0 ^~ inbuffer_data[167];
assign xnor8[168] = 1'b0 ^~ inbuffer_data[168];
assign xnor8[169] = 1'b1 ^~ inbuffer_data[169];
assign xnor8[170] = 1'b1 ^~ inbuffer_data[170];
assign xnor8[171] = 1'b0 ^~ inbuffer_data[171];
assign xnor8[172] = 1'b0 ^~ inbuffer_data[172];
assign xnor8[173] = 1'b1 ^~ inbuffer_data[173];
assign xnor8[174] = 1'b1 ^~ inbuffer_data[174];
assign xnor8[175] = 1'b1 ^~ inbuffer_data[175];
assign xnor8[176] = 1'b1 ^~ inbuffer_data[176];
assign xnor8[177] = 1'b0 ^~ inbuffer_data[177];
assign xnor8[178] = 1'b1 ^~ inbuffer_data[178];
assign xnor8[179] = 1'b0 ^~ inbuffer_data[179];
assign xnor8[180] = 1'b1 ^~ inbuffer_data[180];
assign xnor8[181] = 1'b1 ^~ inbuffer_data[181];
assign xnor8[182] = 1'b1 ^~ inbuffer_data[182];
assign xnor8[183] = 1'b1 ^~ inbuffer_data[183];
assign xnor8[184] = 1'b1 ^~ inbuffer_data[184];
assign xnor8[185] = 1'b1 ^~ inbuffer_data[185];
assign xnor8[186] = 1'b0 ^~ inbuffer_data[186];
assign xnor8[187] = 1'b1 ^~ inbuffer_data[187];
assign xnor8[188] = 1'b1 ^~ inbuffer_data[188];
assign xnor8[189] = 1'b0 ^~ inbuffer_data[189];
assign xnor8[190] = 1'b1 ^~ inbuffer_data[190];
assign xnor8[191] = 1'b1 ^~ inbuffer_data[191];
assign xnor8[192] = 1'b1 ^~ inbuffer_data[192];
assign xnor8[193] = 1'b0 ^~ inbuffer_data[193];
assign xnor8[194] = 1'b1 ^~ inbuffer_data[194];
assign xnor8[195] = 1'b1 ^~ inbuffer_data[195];
assign xnor8[196] = 1'b0 ^~ inbuffer_data[196];
assign xnor8[197] = 1'b0 ^~ inbuffer_data[197];
assign xnor8[198] = 1'b1 ^~ inbuffer_data[198];
assign xnor8[199] = 1'b0 ^~ inbuffer_data[199];
assign xnor8[200] = 1'b0 ^~ inbuffer_data[200];
assign xnor8[201] = 1'b0 ^~ inbuffer_data[201];
assign xnor8[202] = 1'b0 ^~ inbuffer_data[202];
assign xnor8[203] = 1'b0 ^~ inbuffer_data[203];
assign xnor8[204] = 1'b1 ^~ inbuffer_data[204];
assign xnor8[205] = 1'b0 ^~ inbuffer_data[205];
assign xnor8[206] = 1'b1 ^~ inbuffer_data[206];
assign xnor8[207] = 1'b0 ^~ inbuffer_data[207];
assign xnor8[208] = 1'b0 ^~ inbuffer_data[208];
assign xnor8[209] = 1'b0 ^~ inbuffer_data[209];
assign xnor8[210] = 1'b0 ^~ inbuffer_data[210];
assign xnor8[211] = 1'b0 ^~ inbuffer_data[211];
assign xnor8[212] = 1'b0 ^~ inbuffer_data[212];
assign xnor8[213] = 1'b1 ^~ inbuffer_data[213];
assign xnor8[214] = 1'b1 ^~ inbuffer_data[214];
assign xnor8[215] = 1'b1 ^~ inbuffer_data[215];
assign xnor8[216] = 1'b1 ^~ inbuffer_data[216];
assign xnor8[217] = 1'b1 ^~ inbuffer_data[217];
assign xnor8[218] = 1'b0 ^~ inbuffer_data[218];
assign xnor8[219] = 1'b1 ^~ inbuffer_data[219];
assign xnor8[220] = 1'b1 ^~ inbuffer_data[220];
assign xnor8[221] = 1'b1 ^~ inbuffer_data[221];
assign xnor8[222] = 1'b0 ^~ inbuffer_data[222];
assign xnor8[223] = 1'b0 ^~ inbuffer_data[223];
assign xnor8[224] = 1'b1 ^~ inbuffer_data[224];
assign xnor8[225] = 1'b0 ^~ inbuffer_data[225];
assign xnor8[226] = 1'b0 ^~ inbuffer_data[226];
assign xnor8[227] = 1'b1 ^~ inbuffer_data[227];
assign xnor8[228] = 1'b0 ^~ inbuffer_data[228];
assign xnor8[229] = 1'b0 ^~ inbuffer_data[229];
assign xnor8[230] = 1'b1 ^~ inbuffer_data[230];
assign xnor8[231] = 1'b1 ^~ inbuffer_data[231];
assign xnor8[232] = 1'b1 ^~ inbuffer_data[232];
assign xnor8[233] = 1'b1 ^~ inbuffer_data[233];
assign xnor8[234] = 1'b1 ^~ inbuffer_data[234];
assign xnor8[235] = 1'b0 ^~ inbuffer_data[235];
assign xnor8[236] = 1'b1 ^~ inbuffer_data[236];
assign xnor8[237] = 1'b1 ^~ inbuffer_data[237];
assign xnor8[238] = 1'b0 ^~ inbuffer_data[238];
assign xnor8[239] = 1'b0 ^~ inbuffer_data[239];
assign xnor8[240] = 1'b1 ^~ inbuffer_data[240];
assign xnor8[241] = 1'b1 ^~ inbuffer_data[241];
assign xnor8[242] = 1'b1 ^~ inbuffer_data[242];
assign xnor8[243] = 1'b1 ^~ inbuffer_data[243];
assign xnor8[244] = 1'b0 ^~ inbuffer_data[244];
assign xnor8[245] = 1'b1 ^~ inbuffer_data[245];
assign xnor8[246] = 1'b1 ^~ inbuffer_data[246];
assign xnor8[247] = 1'b1 ^~ inbuffer_data[247];
assign xnor8[248] = 1'b1 ^~ inbuffer_data[248];
assign xnor8[249] = 1'b1 ^~ inbuffer_data[249];
assign xnor8[250] = 1'b0 ^~ inbuffer_data[250];
assign xnor8[251] = 1'b1 ^~ inbuffer_data[251];
assign xnor8[252] = 1'b1 ^~ inbuffer_data[252];
assign xnor8[253] = 1'b0 ^~ inbuffer_data[253];
assign xnor8[254] = 1'b1 ^~ inbuffer_data[254];
assign xnor8[255] = 1'b1 ^~ inbuffer_data[255];
assign xnor8[256] = 1'b1 ^~ inbuffer_data[256];
assign xnor8[257] = 1'b1 ^~ inbuffer_data[257];
assign xnor8[258] = 1'b1 ^~ inbuffer_data[258];
assign xnor8[259] = 1'b0 ^~ inbuffer_data[259];
assign xnor8[260] = 1'b1 ^~ inbuffer_data[260];
assign xnor8[261] = 1'b1 ^~ inbuffer_data[261];
assign xnor8[262] = 1'b1 ^~ inbuffer_data[262];
assign xnor8[263] = 1'b1 ^~ inbuffer_data[263];
assign xnor8[264] = 1'b1 ^~ inbuffer_data[264];
assign xnor8[265] = 1'b1 ^~ inbuffer_data[265];
assign xnor8[266] = 1'b0 ^~ inbuffer_data[266];
assign xnor8[267] = 1'b0 ^~ inbuffer_data[267];
assign xnor8[268] = 1'b0 ^~ inbuffer_data[268];
assign xnor8[269] = 1'b1 ^~ inbuffer_data[269];
assign xnor8[270] = 1'b1 ^~ inbuffer_data[270];
assign xnor8[271] = 1'b1 ^~ inbuffer_data[271];
assign xnor8[272] = 1'b1 ^~ inbuffer_data[272];
assign xnor8[273] = 1'b0 ^~ inbuffer_data[273];
assign xnor8[274] = 1'b1 ^~ inbuffer_data[274];
assign xnor8[275] = 1'b1 ^~ inbuffer_data[275];
assign xnor8[276] = 1'b0 ^~ inbuffer_data[276];
assign xnor8[277] = 1'b0 ^~ inbuffer_data[277];
assign xnor8[278] = 1'b1 ^~ inbuffer_data[278];
assign xnor8[279] = 1'b0 ^~ inbuffer_data[279];
assign xnor8[280] = 1'b0 ^~ inbuffer_data[280];
assign xnor8[281] = 1'b0 ^~ inbuffer_data[281];
assign xnor8[282] = 1'b1 ^~ inbuffer_data[282];
assign xnor8[283] = 1'b0 ^~ inbuffer_data[283];
assign xnor8[284] = 1'b1 ^~ inbuffer_data[284];
assign xnor8[285] = 1'b0 ^~ inbuffer_data[285];
assign xnor8[286] = 1'b1 ^~ inbuffer_data[286];
assign xnor8[287] = 1'b1 ^~ inbuffer_data[287];
assign xnor8[288] = 1'b1 ^~ inbuffer_data[288];
assign xnor8[289] = 1'b1 ^~ inbuffer_data[289];
assign xnor8[290] = 1'b1 ^~ inbuffer_data[290];
assign xnor8[291] = 1'b1 ^~ inbuffer_data[291];
assign xnor8[292] = 1'b1 ^~ inbuffer_data[292];
assign xnor8[293] = 1'b1 ^~ inbuffer_data[293];
assign xnor8[294] = 1'b0 ^~ inbuffer_data[294];
assign xnor8[295] = 1'b0 ^~ inbuffer_data[295];
assign xnor8[296] = 1'b0 ^~ inbuffer_data[296];
assign xnor8[297] = 1'b0 ^~ inbuffer_data[297];
assign xnor8[298] = 1'b1 ^~ inbuffer_data[298];
assign xnor8[299] = 1'b1 ^~ inbuffer_data[299];
assign xnor8[300] = 1'b1 ^~ inbuffer_data[300];
assign xnor8[301] = 1'b1 ^~ inbuffer_data[301];
assign xnor8[302] = 1'b1 ^~ inbuffer_data[302];
assign xnor8[303] = 1'b1 ^~ inbuffer_data[303];
assign xnor8[304] = 1'b0 ^~ inbuffer_data[304];
assign xnor8[305] = 1'b0 ^~ inbuffer_data[305];
assign xnor8[306] = 1'b0 ^~ inbuffer_data[306];
assign xnor8[307] = 1'b1 ^~ inbuffer_data[307];
assign xnor8[308] = 1'b0 ^~ inbuffer_data[308];
assign xnor8[309] = 1'b0 ^~ inbuffer_data[309];
assign xnor8[310] = 1'b0 ^~ inbuffer_data[310];
assign xnor8[311] = 1'b0 ^~ inbuffer_data[311];
assign xnor8[312] = 1'b1 ^~ inbuffer_data[312];
assign xnor8[313] = 1'b1 ^~ inbuffer_data[313];
assign xnor8[314] = 1'b1 ^~ inbuffer_data[314];
assign xnor8[315] = 1'b1 ^~ inbuffer_data[315];
assign xnor8[316] = 1'b1 ^~ inbuffer_data[316];
assign xnor8[317] = 1'b1 ^~ inbuffer_data[317];
assign xnor8[318] = 1'b1 ^~ inbuffer_data[318];
assign xnor8[319] = 1'b1 ^~ inbuffer_data[319];
assign xnor8[320] = 1'b1 ^~ inbuffer_data[320];
assign xnor8[321] = 1'b1 ^~ inbuffer_data[321];
assign xnor8[322] = 1'b1 ^~ inbuffer_data[322];
assign xnor8[323] = 1'b1 ^~ inbuffer_data[323];
assign xnor8[324] = 1'b0 ^~ inbuffer_data[324];
assign xnor8[325] = 1'b0 ^~ inbuffer_data[325];
assign xnor8[326] = 1'b0 ^~ inbuffer_data[326];
assign xnor8[327] = 1'b1 ^~ inbuffer_data[327];
assign xnor8[328] = 1'b1 ^~ inbuffer_data[328];
assign xnor8[329] = 1'b1 ^~ inbuffer_data[329];
assign xnor8[330] = 1'b1 ^~ inbuffer_data[330];
assign xnor8[331] = 1'b1 ^~ inbuffer_data[331];
assign xnor8[332] = 1'b1 ^~ inbuffer_data[332];
assign xnor8[333] = 1'b1 ^~ inbuffer_data[333];
assign xnor8[334] = 1'b0 ^~ inbuffer_data[334];
assign xnor8[335] = 1'b0 ^~ inbuffer_data[335];
assign xnor8[336] = 1'b1 ^~ inbuffer_data[336];
assign xnor8[337] = 1'b0 ^~ inbuffer_data[337];
assign xnor8[338] = 1'b1 ^~ inbuffer_data[338];
assign xnor8[339] = 1'b0 ^~ inbuffer_data[339];
assign xnor8[340] = 1'b1 ^~ inbuffer_data[340];
assign xnor8[341] = 1'b1 ^~ inbuffer_data[341];
assign xnor8[342] = 1'b1 ^~ inbuffer_data[342];
assign xnor8[343] = 1'b1 ^~ inbuffer_data[343];
assign xnor8[344] = 1'b1 ^~ inbuffer_data[344];
assign xnor8[345] = 1'b1 ^~ inbuffer_data[345];
assign xnor8[346] = 1'b1 ^~ inbuffer_data[346];
assign xnor8[347] = 1'b1 ^~ inbuffer_data[347];
assign xnor8[348] = 1'b1 ^~ inbuffer_data[348];
assign xnor8[349] = 1'b1 ^~ inbuffer_data[349];
assign xnor8[350] = 1'b1 ^~ inbuffer_data[350];
assign xnor8[351] = 1'b1 ^~ inbuffer_data[351];
assign xnor8[352] = 1'b1 ^~ inbuffer_data[352];
assign xnor8[353] = 1'b0 ^~ inbuffer_data[353];
assign xnor8[354] = 1'b0 ^~ inbuffer_data[354];
assign xnor8[355] = 1'b1 ^~ inbuffer_data[355];
assign xnor8[356] = 1'b1 ^~ inbuffer_data[356];
assign xnor8[357] = 1'b1 ^~ inbuffer_data[357];
assign xnor8[358] = 1'b1 ^~ inbuffer_data[358];
assign xnor8[359] = 1'b1 ^~ inbuffer_data[359];
assign xnor8[360] = 1'b1 ^~ inbuffer_data[360];
assign xnor8[361] = 1'b1 ^~ inbuffer_data[361];
assign xnor8[362] = 1'b1 ^~ inbuffer_data[362];
assign xnor8[363] = 1'b0 ^~ inbuffer_data[363];
assign xnor8[364] = 1'b0 ^~ inbuffer_data[364];
assign xnor8[365] = 1'b1 ^~ inbuffer_data[365];
assign xnor8[366] = 1'b1 ^~ inbuffer_data[366];
assign xnor8[367] = 1'b0 ^~ inbuffer_data[367];
assign xnor8[368] = 1'b0 ^~ inbuffer_data[368];
assign xnor8[369] = 1'b1 ^~ inbuffer_data[369];
assign xnor8[370] = 1'b1 ^~ inbuffer_data[370];
assign xnor8[371] = 1'b1 ^~ inbuffer_data[371];
assign xnor8[372] = 1'b0 ^~ inbuffer_data[372];
assign xnor8[373] = 1'b1 ^~ inbuffer_data[373];
assign xnor8[374] = 1'b0 ^~ inbuffer_data[374];
assign xnor8[375] = 1'b1 ^~ inbuffer_data[375];
assign xnor8[376] = 1'b1 ^~ inbuffer_data[376];
assign xnor8[377] = 1'b1 ^~ inbuffer_data[377];
assign xnor8[378] = 1'b1 ^~ inbuffer_data[378];
assign xnor8[379] = 1'b1 ^~ inbuffer_data[379];
assign xnor8[380] = 1'b1 ^~ inbuffer_data[380];
assign xnor8[381] = 1'b0 ^~ inbuffer_data[381];
assign xnor8[382] = 1'b0 ^~ inbuffer_data[382];
assign xnor8[383] = 1'b0 ^~ inbuffer_data[383];
assign xnor8[384] = 1'b1 ^~ inbuffer_data[384];
assign xnor8[385] = 1'b1 ^~ inbuffer_data[385];
assign xnor8[386] = 1'b1 ^~ inbuffer_data[386];
assign xnor8[387] = 1'b1 ^~ inbuffer_data[387];
assign xnor8[388] = 1'b1 ^~ inbuffer_data[388];
assign xnor8[389] = 1'b0 ^~ inbuffer_data[389];
assign xnor8[390] = 1'b0 ^~ inbuffer_data[390];
assign xnor8[391] = 1'b1 ^~ inbuffer_data[391];
assign xnor8[392] = 1'b0 ^~ inbuffer_data[392];
assign xnor8[393] = 1'b0 ^~ inbuffer_data[393];
assign xnor8[394] = 1'b1 ^~ inbuffer_data[394];
assign xnor8[395] = 1'b1 ^~ inbuffer_data[395];
assign xnor8[396] = 1'b1 ^~ inbuffer_data[396];
assign xnor8[397] = 1'b0 ^~ inbuffer_data[397];
assign xnor8[398] = 1'b0 ^~ inbuffer_data[398];
assign xnor8[399] = 1'b0 ^~ inbuffer_data[399];
assign xnor8[400] = 1'b0 ^~ inbuffer_data[400];
assign xnor8[401] = 1'b0 ^~ inbuffer_data[401];
assign xnor8[402] = 1'b0 ^~ inbuffer_data[402];
assign xnor8[403] = 1'b1 ^~ inbuffer_data[403];
assign xnor8[404] = 1'b1 ^~ inbuffer_data[404];
assign xnor8[405] = 1'b1 ^~ inbuffer_data[405];
assign xnor8[406] = 1'b1 ^~ inbuffer_data[406];
assign xnor8[407] = 1'b1 ^~ inbuffer_data[407];
assign xnor8[408] = 1'b1 ^~ inbuffer_data[408];
assign xnor8[409] = 1'b0 ^~ inbuffer_data[409];
assign xnor8[410] = 1'b0 ^~ inbuffer_data[410];
assign xnor8[411] = 1'b0 ^~ inbuffer_data[411];
assign xnor8[412] = 1'b0 ^~ inbuffer_data[412];
assign xnor8[413] = 1'b1 ^~ inbuffer_data[413];
assign xnor8[414] = 1'b0 ^~ inbuffer_data[414];
assign xnor8[415] = 1'b0 ^~ inbuffer_data[415];
assign xnor8[416] = 1'b0 ^~ inbuffer_data[416];
assign xnor8[417] = 1'b1 ^~ inbuffer_data[417];
assign xnor8[418] = 1'b1 ^~ inbuffer_data[418];
assign xnor8[419] = 1'b1 ^~ inbuffer_data[419];
assign xnor8[420] = 1'b0 ^~ inbuffer_data[420];
assign xnor8[421] = 1'b0 ^~ inbuffer_data[421];
assign xnor8[422] = 1'b0 ^~ inbuffer_data[422];
assign xnor8[423] = 1'b1 ^~ inbuffer_data[423];
assign xnor8[424] = 1'b1 ^~ inbuffer_data[424];
assign xnor8[425] = 1'b0 ^~ inbuffer_data[425];
assign xnor8[426] = 1'b0 ^~ inbuffer_data[426];
assign xnor8[427] = 1'b0 ^~ inbuffer_data[427];
assign xnor8[428] = 1'b0 ^~ inbuffer_data[428];
assign xnor8[429] = 1'b0 ^~ inbuffer_data[429];
assign xnor8[430] = 1'b0 ^~ inbuffer_data[430];
assign xnor8[431] = 1'b1 ^~ inbuffer_data[431];
assign xnor8[432] = 1'b1 ^~ inbuffer_data[432];
assign xnor8[433] = 1'b1 ^~ inbuffer_data[433];
assign xnor8[434] = 1'b1 ^~ inbuffer_data[434];
assign xnor8[435] = 1'b1 ^~ inbuffer_data[435];
assign xnor8[436] = 1'b1 ^~ inbuffer_data[436];
assign xnor8[437] = 1'b1 ^~ inbuffer_data[437];
assign xnor8[438] = 1'b0 ^~ inbuffer_data[438];
assign xnor8[439] = 1'b0 ^~ inbuffer_data[439];
assign xnor8[440] = 1'b1 ^~ inbuffer_data[440];
assign xnor8[441] = 1'b0 ^~ inbuffer_data[441];
assign xnor8[442] = 1'b0 ^~ inbuffer_data[442];
assign xnor8[443] = 1'b0 ^~ inbuffer_data[443];
assign xnor8[444] = 1'b0 ^~ inbuffer_data[444];
assign xnor8[445] = 1'b0 ^~ inbuffer_data[445];
assign xnor8[446] = 1'b0 ^~ inbuffer_data[446];
assign xnor8[447] = 1'b0 ^~ inbuffer_data[447];
assign xnor8[448] = 1'b0 ^~ inbuffer_data[448];
assign xnor8[449] = 1'b1 ^~ inbuffer_data[449];
assign xnor8[450] = 1'b0 ^~ inbuffer_data[450];
assign xnor8[451] = 1'b0 ^~ inbuffer_data[451];
assign xnor8[452] = 1'b0 ^~ inbuffer_data[452];
assign xnor8[453] = 1'b0 ^~ inbuffer_data[453];
assign xnor8[454] = 1'b1 ^~ inbuffer_data[454];
assign xnor8[455] = 1'b0 ^~ inbuffer_data[455];
assign xnor8[456] = 1'b1 ^~ inbuffer_data[456];
assign xnor8[457] = 1'b1 ^~ inbuffer_data[457];
assign xnor8[458] = 1'b0 ^~ inbuffer_data[458];
assign xnor8[459] = 1'b1 ^~ inbuffer_data[459];
assign xnor8[460] = 1'b1 ^~ inbuffer_data[460];
assign xnor8[461] = 1'b1 ^~ inbuffer_data[461];
assign xnor8[462] = 1'b1 ^~ inbuffer_data[462];
assign xnor8[463] = 1'b1 ^~ inbuffer_data[463];
assign xnor8[464] = 1'b0 ^~ inbuffer_data[464];
assign xnor8[465] = 1'b0 ^~ inbuffer_data[465];
assign xnor8[466] = 1'b0 ^~ inbuffer_data[466];
assign xnor8[467] = 1'b0 ^~ inbuffer_data[467];
assign xnor8[468] = 1'b0 ^~ inbuffer_data[468];
assign xnor8[469] = 1'b0 ^~ inbuffer_data[469];
assign xnor8[470] = 1'b0 ^~ inbuffer_data[470];
assign xnor8[471] = 1'b1 ^~ inbuffer_data[471];
assign xnor8[472] = 1'b0 ^~ inbuffer_data[472];
assign xnor8[473] = 1'b1 ^~ inbuffer_data[473];
assign xnor8[474] = 1'b0 ^~ inbuffer_data[474];
assign xnor8[475] = 1'b0 ^~ inbuffer_data[475];
assign xnor8[476] = 1'b0 ^~ inbuffer_data[476];
assign xnor8[477] = 1'b1 ^~ inbuffer_data[477];
assign xnor8[478] = 1'b0 ^~ inbuffer_data[478];
assign xnor8[479] = 1'b1 ^~ inbuffer_data[479];
assign xnor8[480] = 1'b1 ^~ inbuffer_data[480];
assign xnor8[481] = 1'b0 ^~ inbuffer_data[481];
assign xnor8[482] = 1'b0 ^~ inbuffer_data[482];
assign xnor8[483] = 1'b1 ^~ inbuffer_data[483];
assign xnor8[484] = 1'b1 ^~ inbuffer_data[484];
assign xnor8[485] = 1'b1 ^~ inbuffer_data[485];
assign xnor8[486] = 1'b1 ^~ inbuffer_data[486];
assign xnor8[487] = 1'b1 ^~ inbuffer_data[487];
assign xnor8[488] = 1'b1 ^~ inbuffer_data[488];
assign xnor8[489] = 1'b1 ^~ inbuffer_data[489];
assign xnor8[490] = 1'b1 ^~ inbuffer_data[490];
assign xnor8[491] = 1'b0 ^~ inbuffer_data[491];
assign xnor8[492] = 1'b1 ^~ inbuffer_data[492];
assign xnor8[493] = 1'b0 ^~ inbuffer_data[493];
assign xnor8[494] = 1'b0 ^~ inbuffer_data[494];
assign xnor8[495] = 1'b0 ^~ inbuffer_data[495];
assign xnor8[496] = 1'b0 ^~ inbuffer_data[496];
assign xnor8[497] = 1'b0 ^~ inbuffer_data[497];
assign xnor8[498] = 1'b0 ^~ inbuffer_data[498];
assign xnor8[499] = 1'b1 ^~ inbuffer_data[499];
assign xnor8[500] = 1'b1 ^~ inbuffer_data[500];
assign xnor8[501] = 1'b0 ^~ inbuffer_data[501];
assign xnor8[502] = 1'b0 ^~ inbuffer_data[502];
assign xnor8[503] = 1'b0 ^~ inbuffer_data[503];
assign xnor8[504] = 1'b1 ^~ inbuffer_data[504];
assign xnor8[505] = 1'b0 ^~ inbuffer_data[505];
assign xnor8[506] = 1'b1 ^~ inbuffer_data[506];
assign xnor8[507] = 1'b0 ^~ inbuffer_data[507];
assign xnor8[508] = 1'b0 ^~ inbuffer_data[508];
assign xnor8[509] = 1'b1 ^~ inbuffer_data[509];
assign xnor8[510] = 1'b1 ^~ inbuffer_data[510];
assign xnor8[511] = 1'b1 ^~ inbuffer_data[511];
assign xnor8[512] = 1'b1 ^~ inbuffer_data[512];
assign xnor8[513] = 1'b1 ^~ inbuffer_data[513];
assign xnor8[514] = 1'b1 ^~ inbuffer_data[514];
assign xnor8[515] = 1'b1 ^~ inbuffer_data[515];
assign xnor8[516] = 1'b1 ^~ inbuffer_data[516];
assign xnor8[517] = 1'b1 ^~ inbuffer_data[517];
assign xnor8[518] = 1'b0 ^~ inbuffer_data[518];
assign xnor8[519] = 1'b0 ^~ inbuffer_data[519];
assign xnor8[520] = 1'b1 ^~ inbuffer_data[520];
assign xnor8[521] = 1'b0 ^~ inbuffer_data[521];
assign xnor8[522] = 1'b0 ^~ inbuffer_data[522];
assign xnor8[523] = 1'b1 ^~ inbuffer_data[523];
assign xnor8[524] = 1'b0 ^~ inbuffer_data[524];
assign xnor8[525] = 1'b0 ^~ inbuffer_data[525];
assign xnor8[526] = 1'b1 ^~ inbuffer_data[526];
assign xnor8[527] = 1'b0 ^~ inbuffer_data[527];
assign xnor8[528] = 1'b0 ^~ inbuffer_data[528];
assign xnor8[529] = 1'b0 ^~ inbuffer_data[529];
assign xnor8[530] = 1'b0 ^~ inbuffer_data[530];
assign xnor8[531] = 1'b0 ^~ inbuffer_data[531];
assign xnor8[532] = 1'b0 ^~ inbuffer_data[532];
assign xnor8[533] = 1'b1 ^~ inbuffer_data[533];
assign xnor8[534] = 1'b0 ^~ inbuffer_data[534];
assign xnor8[535] = 1'b0 ^~ inbuffer_data[535];
assign xnor8[536] = 1'b0 ^~ inbuffer_data[536];
assign xnor8[537] = 1'b1 ^~ inbuffer_data[537];
assign xnor8[538] = 1'b0 ^~ inbuffer_data[538];
assign xnor8[539] = 1'b1 ^~ inbuffer_data[539];
assign xnor8[540] = 1'b1 ^~ inbuffer_data[540];
assign xnor8[541] = 1'b1 ^~ inbuffer_data[541];
assign xnor8[542] = 1'b1 ^~ inbuffer_data[542];
assign xnor8[543] = 1'b0 ^~ inbuffer_data[543];
assign xnor8[544] = 1'b0 ^~ inbuffer_data[544];
assign xnor8[545] = 1'b0 ^~ inbuffer_data[545];
assign xnor8[546] = 1'b0 ^~ inbuffer_data[546];
assign xnor8[547] = 1'b1 ^~ inbuffer_data[547];
assign xnor8[548] = 1'b0 ^~ inbuffer_data[548];
assign xnor8[549] = 1'b0 ^~ inbuffer_data[549];
assign xnor8[550] = 1'b1 ^~ inbuffer_data[550];
assign xnor8[551] = 1'b1 ^~ inbuffer_data[551];
assign xnor8[552] = 1'b0 ^~ inbuffer_data[552];
assign xnor8[553] = 1'b1 ^~ inbuffer_data[553];
assign xnor8[554] = 1'b1 ^~ inbuffer_data[554];
assign xnor8[555] = 1'b1 ^~ inbuffer_data[555];
assign xnor8[556] = 1'b0 ^~ inbuffer_data[556];
assign xnor8[557] = 1'b1 ^~ inbuffer_data[557];
assign xnor8[558] = 1'b0 ^~ inbuffer_data[558];
assign xnor8[559] = 1'b0 ^~ inbuffer_data[559];
assign xnor8[560] = 1'b1 ^~ inbuffer_data[560];
assign xnor8[561] = 1'b0 ^~ inbuffer_data[561];
assign xnor8[562] = 1'b1 ^~ inbuffer_data[562];
assign xnor8[563] = 1'b1 ^~ inbuffer_data[563];
assign xnor8[564] = 1'b0 ^~ inbuffer_data[564];
assign xnor8[565] = 1'b1 ^~ inbuffer_data[565];
assign xnor8[566] = 1'b1 ^~ inbuffer_data[566];
assign xnor8[567] = 1'b1 ^~ inbuffer_data[567];
assign xnor8[568] = 1'b0 ^~ inbuffer_data[568];
assign xnor8[569] = 1'b1 ^~ inbuffer_data[569];
assign xnor8[570] = 1'b1 ^~ inbuffer_data[570];
assign xnor8[571] = 1'b0 ^~ inbuffer_data[571];
assign xnor8[572] = 1'b0 ^~ inbuffer_data[572];
assign xnor8[573] = 1'b1 ^~ inbuffer_data[573];
assign xnor8[574] = 1'b0 ^~ inbuffer_data[574];
assign xnor8[575] = 1'b1 ^~ inbuffer_data[575];
assign xnor8[576] = 1'b0 ^~ inbuffer_data[576];
assign xnor8[577] = 1'b0 ^~ inbuffer_data[577];
assign xnor8[578] = 1'b1 ^~ inbuffer_data[578];
assign xnor8[579] = 1'b1 ^~ inbuffer_data[579];
assign xnor8[580] = 1'b1 ^~ inbuffer_data[580];
assign xnor8[581] = 1'b1 ^~ inbuffer_data[581];
assign xnor8[582] = 1'b1 ^~ inbuffer_data[582];
assign xnor8[583] = 1'b0 ^~ inbuffer_data[583];
assign xnor8[584] = 1'b0 ^~ inbuffer_data[584];
assign xnor8[585] = 1'b0 ^~ inbuffer_data[585];
assign xnor8[586] = 1'b0 ^~ inbuffer_data[586];
assign xnor8[587] = 1'b1 ^~ inbuffer_data[587];
assign xnor8[588] = 1'b1 ^~ inbuffer_data[588];
assign xnor8[589] = 1'b0 ^~ inbuffer_data[589];
assign xnor8[590] = 1'b1 ^~ inbuffer_data[590];
assign xnor8[591] = 1'b0 ^~ inbuffer_data[591];
assign xnor8[592] = 1'b0 ^~ inbuffer_data[592];
assign xnor8[593] = 1'b1 ^~ inbuffer_data[593];
assign xnor8[594] = 1'b1 ^~ inbuffer_data[594];
assign xnor8[595] = 1'b1 ^~ inbuffer_data[595];
assign xnor8[596] = 1'b0 ^~ inbuffer_data[596];
assign xnor8[597] = 1'b1 ^~ inbuffer_data[597];
assign xnor8[598] = 1'b1 ^~ inbuffer_data[598];
assign xnor8[599] = 1'b0 ^~ inbuffer_data[599];
assign xnor8[600] = 1'b0 ^~ inbuffer_data[600];
assign xnor8[601] = 1'b0 ^~ inbuffer_data[601];
assign xnor8[602] = 1'b0 ^~ inbuffer_data[602];
assign xnor8[603] = 1'b0 ^~ inbuffer_data[603];
assign xnor8[604] = 1'b0 ^~ inbuffer_data[604];
assign xnor8[605] = 1'b0 ^~ inbuffer_data[605];
assign xnor8[606] = 1'b1 ^~ inbuffer_data[606];
assign xnor8[607] = 1'b0 ^~ inbuffer_data[607];
assign xnor8[608] = 1'b1 ^~ inbuffer_data[608];
assign xnor8[609] = 1'b1 ^~ inbuffer_data[609];
assign xnor8[610] = 1'b1 ^~ inbuffer_data[610];
assign xnor8[611] = 1'b0 ^~ inbuffer_data[611];
assign xnor8[612] = 1'b0 ^~ inbuffer_data[612];
assign xnor8[613] = 1'b0 ^~ inbuffer_data[613];
assign xnor8[614] = 1'b1 ^~ inbuffer_data[614];
assign xnor8[615] = 1'b1 ^~ inbuffer_data[615];
assign xnor8[616] = 1'b1 ^~ inbuffer_data[616];
assign xnor8[617] = 1'b1 ^~ inbuffer_data[617];
assign xnor8[618] = 1'b0 ^~ inbuffer_data[618];
assign xnor8[619] = 1'b1 ^~ inbuffer_data[619];
assign xnor8[620] = 1'b0 ^~ inbuffer_data[620];
assign xnor8[621] = 1'b0 ^~ inbuffer_data[621];
assign xnor8[622] = 1'b0 ^~ inbuffer_data[622];
assign xnor8[623] = 1'b1 ^~ inbuffer_data[623];
assign xnor8[624] = 1'b1 ^~ inbuffer_data[624];
assign xnor8[625] = 1'b0 ^~ inbuffer_data[625];
assign xnor8[626] = 1'b0 ^~ inbuffer_data[626];
assign xnor8[627] = 1'b0 ^~ inbuffer_data[627];
assign xnor8[628] = 1'b1 ^~ inbuffer_data[628];
assign xnor8[629] = 1'b1 ^~ inbuffer_data[629];
assign xnor8[630] = 1'b1 ^~ inbuffer_data[630];
assign xnor8[631] = 1'b1 ^~ inbuffer_data[631];
assign xnor8[632] = 1'b1 ^~ inbuffer_data[632];
assign xnor8[633] = 1'b0 ^~ inbuffer_data[633];
assign xnor8[634] = 1'b1 ^~ inbuffer_data[634];
assign xnor8[635] = 1'b1 ^~ inbuffer_data[635];
assign xnor8[636] = 1'b1 ^~ inbuffer_data[636];
assign xnor8[637] = 1'b1 ^~ inbuffer_data[637];
assign xnor8[638] = 1'b0 ^~ inbuffer_data[638];
assign xnor8[639] = 1'b1 ^~ inbuffer_data[639];
assign xnor8[640] = 1'b0 ^~ inbuffer_data[640];
assign xnor8[641] = 1'b0 ^~ inbuffer_data[641];
assign xnor8[642] = 1'b0 ^~ inbuffer_data[642];
assign xnor8[643] = 1'b0 ^~ inbuffer_data[643];
assign xnor8[644] = 1'b0 ^~ inbuffer_data[644];
assign xnor8[645] = 1'b1 ^~ inbuffer_data[645];
assign xnor8[646] = 1'b1 ^~ inbuffer_data[646];
assign xnor8[647] = 1'b0 ^~ inbuffer_data[647];
assign xnor8[648] = 1'b1 ^~ inbuffer_data[648];
assign xnor8[649] = 1'b0 ^~ inbuffer_data[649];
assign xnor8[650] = 1'b0 ^~ inbuffer_data[650];
assign xnor8[651] = 1'b0 ^~ inbuffer_data[651];
assign xnor8[652] = 1'b1 ^~ inbuffer_data[652];
assign xnor8[653] = 1'b1 ^~ inbuffer_data[653];
assign xnor8[654] = 1'b1 ^~ inbuffer_data[654];
assign xnor8[655] = 1'b0 ^~ inbuffer_data[655];
assign xnor8[656] = 1'b1 ^~ inbuffer_data[656];
assign xnor8[657] = 1'b1 ^~ inbuffer_data[657];
assign xnor8[658] = 1'b1 ^~ inbuffer_data[658];
assign xnor8[659] = 1'b1 ^~ inbuffer_data[659];
assign xnor8[660] = 1'b1 ^~ inbuffer_data[660];
assign xnor8[661] = 1'b0 ^~ inbuffer_data[661];
assign xnor8[662] = 1'b1 ^~ inbuffer_data[662];
assign xnor8[663] = 1'b1 ^~ inbuffer_data[663];
assign xnor8[664] = 1'b1 ^~ inbuffer_data[664];
assign xnor8[665] = 1'b0 ^~ inbuffer_data[665];
assign xnor8[666] = 1'b0 ^~ inbuffer_data[666];
assign xnor8[667] = 1'b0 ^~ inbuffer_data[667];
assign xnor8[668] = 1'b0 ^~ inbuffer_data[668];
assign xnor8[669] = 1'b0 ^~ inbuffer_data[669];
assign xnor8[670] = 1'b0 ^~ inbuffer_data[670];
assign xnor8[671] = 1'b0 ^~ inbuffer_data[671];
assign xnor8[672] = 1'b0 ^~ inbuffer_data[672];
assign xnor8[673] = 1'b0 ^~ inbuffer_data[673];
assign xnor8[674] = 1'b1 ^~ inbuffer_data[674];
assign xnor8[675] = 1'b1 ^~ inbuffer_data[675];
assign xnor8[676] = 1'b0 ^~ inbuffer_data[676];
assign xnor8[677] = 1'b0 ^~ inbuffer_data[677];
assign xnor8[678] = 1'b0 ^~ inbuffer_data[678];
assign xnor8[679] = 1'b0 ^~ inbuffer_data[679];
assign xnor8[680] = 1'b0 ^~ inbuffer_data[680];
assign xnor8[681] = 1'b1 ^~ inbuffer_data[681];
assign xnor8[682] = 1'b1 ^~ inbuffer_data[682];
assign xnor8[683] = 1'b1 ^~ inbuffer_data[683];
assign xnor8[684] = 1'b1 ^~ inbuffer_data[684];
assign xnor8[685] = 1'b1 ^~ inbuffer_data[685];
assign xnor8[686] = 1'b1 ^~ inbuffer_data[686];
assign xnor8[687] = 1'b1 ^~ inbuffer_data[687];
assign xnor8[688] = 1'b1 ^~ inbuffer_data[688];
assign xnor8[689] = 1'b1 ^~ inbuffer_data[689];
assign xnor8[690] = 1'b1 ^~ inbuffer_data[690];
assign xnor8[691] = 1'b1 ^~ inbuffer_data[691];
assign xnor8[692] = 1'b1 ^~ inbuffer_data[692];
assign xnor8[693] = 1'b0 ^~ inbuffer_data[693];
assign xnor8[694] = 1'b1 ^~ inbuffer_data[694];
assign xnor8[695] = 1'b0 ^~ inbuffer_data[695];
assign xnor8[696] = 1'b1 ^~ inbuffer_data[696];
assign xnor8[697] = 1'b1 ^~ inbuffer_data[697];
assign xnor8[698] = 1'b1 ^~ inbuffer_data[698];
assign xnor8[699] = 1'b0 ^~ inbuffer_data[699];
assign xnor8[700] = 1'b1 ^~ inbuffer_data[700];
assign xnor8[701] = 1'b1 ^~ inbuffer_data[701];
assign xnor8[702] = 1'b1 ^~ inbuffer_data[702];
assign xnor8[703] = 1'b1 ^~ inbuffer_data[703];
assign xnor8[704] = 1'b1 ^~ inbuffer_data[704];
assign xnor8[705] = 1'b0 ^~ inbuffer_data[705];
assign xnor8[706] = 1'b1 ^~ inbuffer_data[706];
assign xnor8[707] = 1'b0 ^~ inbuffer_data[707];
assign xnor8[708] = 1'b0 ^~ inbuffer_data[708];
assign xnor8[709] = 1'b0 ^~ inbuffer_data[709];
assign xnor8[710] = 1'b0 ^~ inbuffer_data[710];
assign xnor8[711] = 1'b0 ^~ inbuffer_data[711];
assign xnor8[712] = 1'b0 ^~ inbuffer_data[712];
assign xnor8[713] = 1'b1 ^~ inbuffer_data[713];
assign xnor8[714] = 1'b1 ^~ inbuffer_data[714];
assign xnor8[715] = 1'b1 ^~ inbuffer_data[715];
assign xnor8[716] = 1'b1 ^~ inbuffer_data[716];
assign xnor8[717] = 1'b1 ^~ inbuffer_data[717];
assign xnor8[718] = 1'b1 ^~ inbuffer_data[718];
assign xnor8[719] = 1'b0 ^~ inbuffer_data[719];
assign xnor8[720] = 1'b1 ^~ inbuffer_data[720];
assign xnor8[721] = 1'b0 ^~ inbuffer_data[721];
assign xnor8[722] = 1'b1 ^~ inbuffer_data[722];
assign xnor8[723] = 1'b0 ^~ inbuffer_data[723];
assign xnor8[724] = 1'b0 ^~ inbuffer_data[724];
assign xnor8[725] = 1'b0 ^~ inbuffer_data[725];
assign xnor8[726] = 1'b0 ^~ inbuffer_data[726];
assign xnor8[727] = 1'b1 ^~ inbuffer_data[727];
assign xnor8[728] = 1'b1 ^~ inbuffer_data[728];
assign xnor8[729] = 1'b0 ^~ inbuffer_data[729];
assign xnor8[730] = 1'b1 ^~ inbuffer_data[730];
assign xnor8[731] = 1'b0 ^~ inbuffer_data[731];
assign xnor8[732] = 1'b0 ^~ inbuffer_data[732];
assign xnor8[733] = 1'b1 ^~ inbuffer_data[733];
assign xnor8[734] = 1'b0 ^~ inbuffer_data[734];
assign xnor8[735] = 1'b1 ^~ inbuffer_data[735];
assign xnor8[736] = 1'b0 ^~ inbuffer_data[736];
assign xnor8[737] = 1'b0 ^~ inbuffer_data[737];
assign xnor8[738] = 1'b0 ^~ inbuffer_data[738];
assign xnor8[739] = 1'b0 ^~ inbuffer_data[739];
assign xnor8[740] = 1'b0 ^~ inbuffer_data[740];
assign xnor8[741] = 1'b0 ^~ inbuffer_data[741];
assign xnor8[742] = 1'b0 ^~ inbuffer_data[742];
assign xnor8[743] = 1'b0 ^~ inbuffer_data[743];
assign xnor8[744] = 1'b1 ^~ inbuffer_data[744];
assign xnor8[745] = 1'b1 ^~ inbuffer_data[745];
assign xnor8[746] = 1'b0 ^~ inbuffer_data[746];
assign xnor8[747] = 1'b1 ^~ inbuffer_data[747];
assign xnor8[748] = 1'b0 ^~ inbuffer_data[748];
assign xnor8[749] = 1'b1 ^~ inbuffer_data[749];
assign xnor8[750] = 1'b0 ^~ inbuffer_data[750];
assign xnor8[751] = 1'b1 ^~ inbuffer_data[751];
assign xnor8[752] = 1'b1 ^~ inbuffer_data[752];
assign xnor8[753] = 1'b0 ^~ inbuffer_data[753];
assign xnor8[754] = 1'b1 ^~ inbuffer_data[754];
assign xnor8[755] = 1'b0 ^~ inbuffer_data[755];
assign xnor8[756] = 1'b0 ^~ inbuffer_data[756];
assign xnor8[757] = 1'b0 ^~ inbuffer_data[757];
assign xnor8[758] = 1'b1 ^~ inbuffer_data[758];
assign xnor8[759] = 1'b1 ^~ inbuffer_data[759];
assign xnor8[760] = 1'b0 ^~ inbuffer_data[760];
assign xnor8[761] = 1'b0 ^~ inbuffer_data[761];
assign xnor8[762] = 1'b1 ^~ inbuffer_data[762];
assign xnor8[763] = 1'b1 ^~ inbuffer_data[763];
assign xnor8[764] = 1'b0 ^~ inbuffer_data[764];
assign xnor8[765] = 1'b0 ^~ inbuffer_data[765];
assign xnor8[766] = 1'b0 ^~ inbuffer_data[766];
assign xnor8[767] = 1'b1 ^~ inbuffer_data[767];
assign xnor8[768] = 1'b1 ^~ inbuffer_data[768];
assign xnor8[769] = 1'b0 ^~ inbuffer_data[769];
assign xnor8[770] = 1'b0 ^~ inbuffer_data[770];
assign xnor8[771] = 1'b1 ^~ inbuffer_data[771];
assign xnor8[772] = 1'b0 ^~ inbuffer_data[772];
assign xnor8[773] = 1'b1 ^~ inbuffer_data[773];
assign xnor8[774] = 1'b0 ^~ inbuffer_data[774];
assign xnor8[775] = 1'b1 ^~ inbuffer_data[775];
assign xnor8[776] = 1'b0 ^~ inbuffer_data[776];
assign xnor8[777] = 1'b0 ^~ inbuffer_data[777];
assign xnor8[778] = 1'b0 ^~ inbuffer_data[778];
assign xnor8[779] = 1'b0 ^~ inbuffer_data[779];
assign xnor8[780] = 1'b0 ^~ inbuffer_data[780];
assign xnor8[781] = 1'b1 ^~ inbuffer_data[781];
assign xnor8[782] = 1'b0 ^~ inbuffer_data[782];
assign xnor8[783] = 1'b1 ^~ inbuffer_data[783];
assign xnor9[0] = 1'b0 ^~ inbuffer_data[0];
assign xnor9[1] = 1'b1 ^~ inbuffer_data[1];
assign xnor9[2] = 1'b0 ^~ inbuffer_data[2];
assign xnor9[3] = 1'b0 ^~ inbuffer_data[3];
assign xnor9[4] = 1'b1 ^~ inbuffer_data[4];
assign xnor9[5] = 1'b1 ^~ inbuffer_data[5];
assign xnor9[6] = 1'b0 ^~ inbuffer_data[6];
assign xnor9[7] = 1'b1 ^~ inbuffer_data[7];
assign xnor9[8] = 1'b1 ^~ inbuffer_data[8];
assign xnor9[9] = 1'b0 ^~ inbuffer_data[9];
assign xnor9[10] = 1'b0 ^~ inbuffer_data[10];
assign xnor9[11] = 1'b0 ^~ inbuffer_data[11];
assign xnor9[12] = 1'b1 ^~ inbuffer_data[12];
assign xnor9[13] = 1'b0 ^~ inbuffer_data[13];
assign xnor9[14] = 1'b1 ^~ inbuffer_data[14];
assign xnor9[15] = 1'b1 ^~ inbuffer_data[15];
assign xnor9[16] = 1'b0 ^~ inbuffer_data[16];
assign xnor9[17] = 1'b0 ^~ inbuffer_data[17];
assign xnor9[18] = 1'b1 ^~ inbuffer_data[18];
assign xnor9[19] = 1'b0 ^~ inbuffer_data[19];
assign xnor9[20] = 1'b1 ^~ inbuffer_data[20];
assign xnor9[21] = 1'b1 ^~ inbuffer_data[21];
assign xnor9[22] = 1'b0 ^~ inbuffer_data[22];
assign xnor9[23] = 1'b1 ^~ inbuffer_data[23];
assign xnor9[24] = 1'b0 ^~ inbuffer_data[24];
assign xnor9[25] = 1'b0 ^~ inbuffer_data[25];
assign xnor9[26] = 1'b1 ^~ inbuffer_data[26];
assign xnor9[27] = 1'b0 ^~ inbuffer_data[27];
assign xnor9[28] = 1'b1 ^~ inbuffer_data[28];
assign xnor9[29] = 1'b0 ^~ inbuffer_data[29];
assign xnor9[30] = 1'b0 ^~ inbuffer_data[30];
assign xnor9[31] = 1'b1 ^~ inbuffer_data[31];
assign xnor9[32] = 1'b1 ^~ inbuffer_data[32];
assign xnor9[33] = 1'b1 ^~ inbuffer_data[33];
assign xnor9[34] = 1'b1 ^~ inbuffer_data[34];
assign xnor9[35] = 1'b0 ^~ inbuffer_data[35];
assign xnor9[36] = 1'b1 ^~ inbuffer_data[36];
assign xnor9[37] = 1'b0 ^~ inbuffer_data[37];
assign xnor9[38] = 1'b1 ^~ inbuffer_data[38];
assign xnor9[39] = 1'b1 ^~ inbuffer_data[39];
assign xnor9[40] = 1'b1 ^~ inbuffer_data[40];
assign xnor9[41] = 1'b1 ^~ inbuffer_data[41];
assign xnor9[42] = 1'b1 ^~ inbuffer_data[42];
assign xnor9[43] = 1'b0 ^~ inbuffer_data[43];
assign xnor9[44] = 1'b1 ^~ inbuffer_data[44];
assign xnor9[45] = 1'b1 ^~ inbuffer_data[45];
assign xnor9[46] = 1'b1 ^~ inbuffer_data[46];
assign xnor9[47] = 1'b1 ^~ inbuffer_data[47];
assign xnor9[48] = 1'b0 ^~ inbuffer_data[48];
assign xnor9[49] = 1'b0 ^~ inbuffer_data[49];
assign xnor9[50] = 1'b0 ^~ inbuffer_data[50];
assign xnor9[51] = 1'b0 ^~ inbuffer_data[51];
assign xnor9[52] = 1'b1 ^~ inbuffer_data[52];
assign xnor9[53] = 1'b1 ^~ inbuffer_data[53];
assign xnor9[54] = 1'b0 ^~ inbuffer_data[54];
assign xnor9[55] = 1'b1 ^~ inbuffer_data[55];
assign xnor9[56] = 1'b0 ^~ inbuffer_data[56];
assign xnor9[57] = 1'b1 ^~ inbuffer_data[57];
assign xnor9[58] = 1'b1 ^~ inbuffer_data[58];
assign xnor9[59] = 1'b1 ^~ inbuffer_data[59];
assign xnor9[60] = 1'b0 ^~ inbuffer_data[60];
assign xnor9[61] = 1'b0 ^~ inbuffer_data[61];
assign xnor9[62] = 1'b1 ^~ inbuffer_data[62];
assign xnor9[63] = 1'b0 ^~ inbuffer_data[63];
assign xnor9[64] = 1'b0 ^~ inbuffer_data[64];
assign xnor9[65] = 1'b0 ^~ inbuffer_data[65];
assign xnor9[66] = 1'b0 ^~ inbuffer_data[66];
assign xnor9[67] = 1'b1 ^~ inbuffer_data[67];
assign xnor9[68] = 1'b0 ^~ inbuffer_data[68];
assign xnor9[69] = 1'b0 ^~ inbuffer_data[69];
assign xnor9[70] = 1'b0 ^~ inbuffer_data[70];
assign xnor9[71] = 1'b0 ^~ inbuffer_data[71];
assign xnor9[72] = 1'b0 ^~ inbuffer_data[72];
assign xnor9[73] = 1'b0 ^~ inbuffer_data[73];
assign xnor9[74] = 1'b0 ^~ inbuffer_data[74];
assign xnor9[75] = 1'b1 ^~ inbuffer_data[75];
assign xnor9[76] = 1'b0 ^~ inbuffer_data[76];
assign xnor9[77] = 1'b0 ^~ inbuffer_data[77];
assign xnor9[78] = 1'b0 ^~ inbuffer_data[78];
assign xnor9[79] = 1'b0 ^~ inbuffer_data[79];
assign xnor9[80] = 1'b1 ^~ inbuffer_data[80];
assign xnor9[81] = 1'b1 ^~ inbuffer_data[81];
assign xnor9[82] = 1'b1 ^~ inbuffer_data[82];
assign xnor9[83] = 1'b0 ^~ inbuffer_data[83];
assign xnor9[84] = 1'b1 ^~ inbuffer_data[84];
assign xnor9[85] = 1'b1 ^~ inbuffer_data[85];
assign xnor9[86] = 1'b0 ^~ inbuffer_data[86];
assign xnor9[87] = 1'b0 ^~ inbuffer_data[87];
assign xnor9[88] = 1'b0 ^~ inbuffer_data[88];
assign xnor9[89] = 1'b0 ^~ inbuffer_data[89];
assign xnor9[90] = 1'b0 ^~ inbuffer_data[90];
assign xnor9[91] = 1'b0 ^~ inbuffer_data[91];
assign xnor9[92] = 1'b0 ^~ inbuffer_data[92];
assign xnor9[93] = 1'b1 ^~ inbuffer_data[93];
assign xnor9[94] = 1'b1 ^~ inbuffer_data[94];
assign xnor9[95] = 1'b1 ^~ inbuffer_data[95];
assign xnor9[96] = 1'b0 ^~ inbuffer_data[96];
assign xnor9[97] = 1'b1 ^~ inbuffer_data[97];
assign xnor9[98] = 1'b1 ^~ inbuffer_data[98];
assign xnor9[99] = 1'b0 ^~ inbuffer_data[99];
assign xnor9[100] = 1'b0 ^~ inbuffer_data[100];
assign xnor9[101] = 1'b0 ^~ inbuffer_data[101];
assign xnor9[102] = 1'b1 ^~ inbuffer_data[102];
assign xnor9[103] = 1'b1 ^~ inbuffer_data[103];
assign xnor9[104] = 1'b0 ^~ inbuffer_data[104];
assign xnor9[105] = 1'b0 ^~ inbuffer_data[105];
assign xnor9[106] = 1'b0 ^~ inbuffer_data[106];
assign xnor9[107] = 1'b1 ^~ inbuffer_data[107];
assign xnor9[108] = 1'b0 ^~ inbuffer_data[108];
assign xnor9[109] = 1'b0 ^~ inbuffer_data[109];
assign xnor9[110] = 1'b1 ^~ inbuffer_data[110];
assign xnor9[111] = 1'b1 ^~ inbuffer_data[111];
assign xnor9[112] = 1'b0 ^~ inbuffer_data[112];
assign xnor9[113] = 1'b1 ^~ inbuffer_data[113];
assign xnor9[114] = 1'b1 ^~ inbuffer_data[114];
assign xnor9[115] = 1'b0 ^~ inbuffer_data[115];
assign xnor9[116] = 1'b1 ^~ inbuffer_data[116];
assign xnor9[117] = 1'b0 ^~ inbuffer_data[117];
assign xnor9[118] = 1'b1 ^~ inbuffer_data[118];
assign xnor9[119] = 1'b0 ^~ inbuffer_data[119];
assign xnor9[120] = 1'b0 ^~ inbuffer_data[120];
assign xnor9[121] = 1'b0 ^~ inbuffer_data[121];
assign xnor9[122] = 1'b0 ^~ inbuffer_data[122];
assign xnor9[123] = 1'b0 ^~ inbuffer_data[123];
assign xnor9[124] = 1'b0 ^~ inbuffer_data[124];
assign xnor9[125] = 1'b0 ^~ inbuffer_data[125];
assign xnor9[126] = 1'b0 ^~ inbuffer_data[126];
assign xnor9[127] = 1'b0 ^~ inbuffer_data[127];
assign xnor9[128] = 1'b0 ^~ inbuffer_data[128];
assign xnor9[129] = 1'b0 ^~ inbuffer_data[129];
assign xnor9[130] = 1'b0 ^~ inbuffer_data[130];
assign xnor9[131] = 1'b0 ^~ inbuffer_data[131];
assign xnor9[132] = 1'b0 ^~ inbuffer_data[132];
assign xnor9[133] = 1'b0 ^~ inbuffer_data[133];
assign xnor9[134] = 1'b1 ^~ inbuffer_data[134];
assign xnor9[135] = 1'b1 ^~ inbuffer_data[135];
assign xnor9[136] = 1'b1 ^~ inbuffer_data[136];
assign xnor9[137] = 1'b1 ^~ inbuffer_data[137];
assign xnor9[138] = 1'b0 ^~ inbuffer_data[138];
assign xnor9[139] = 1'b1 ^~ inbuffer_data[139];
assign xnor9[140] = 1'b1 ^~ inbuffer_data[140];
assign xnor9[141] = 1'b1 ^~ inbuffer_data[141];
assign xnor9[142] = 1'b1 ^~ inbuffer_data[142];
assign xnor9[143] = 1'b0 ^~ inbuffer_data[143];
assign xnor9[144] = 1'b1 ^~ inbuffer_data[144];
assign xnor9[145] = 1'b1 ^~ inbuffer_data[145];
assign xnor9[146] = 1'b0 ^~ inbuffer_data[146];
assign xnor9[147] = 1'b1 ^~ inbuffer_data[147];
assign xnor9[148] = 1'b1 ^~ inbuffer_data[148];
assign xnor9[149] = 1'b0 ^~ inbuffer_data[149];
assign xnor9[150] = 1'b0 ^~ inbuffer_data[150];
assign xnor9[151] = 1'b1 ^~ inbuffer_data[151];
assign xnor9[152] = 1'b0 ^~ inbuffer_data[152];
assign xnor9[153] = 1'b1 ^~ inbuffer_data[153];
assign xnor9[154] = 1'b0 ^~ inbuffer_data[154];
assign xnor9[155] = 1'b0 ^~ inbuffer_data[155];
assign xnor9[156] = 1'b0 ^~ inbuffer_data[156];
assign xnor9[157] = 1'b0 ^~ inbuffer_data[157];
assign xnor9[158] = 1'b0 ^~ inbuffer_data[158];
assign xnor9[159] = 1'b0 ^~ inbuffer_data[159];
assign xnor9[160] = 1'b0 ^~ inbuffer_data[160];
assign xnor9[161] = 1'b0 ^~ inbuffer_data[161];
assign xnor9[162] = 1'b0 ^~ inbuffer_data[162];
assign xnor9[163] = 1'b1 ^~ inbuffer_data[163];
assign xnor9[164] = 1'b1 ^~ inbuffer_data[164];
assign xnor9[165] = 1'b1 ^~ inbuffer_data[165];
assign xnor9[166] = 1'b1 ^~ inbuffer_data[166];
assign xnor9[167] = 1'b1 ^~ inbuffer_data[167];
assign xnor9[168] = 1'b0 ^~ inbuffer_data[168];
assign xnor9[169] = 1'b1 ^~ inbuffer_data[169];
assign xnor9[170] = 1'b1 ^~ inbuffer_data[170];
assign xnor9[171] = 1'b0 ^~ inbuffer_data[171];
assign xnor9[172] = 1'b1 ^~ inbuffer_data[172];
assign xnor9[173] = 1'b1 ^~ inbuffer_data[173];
assign xnor9[174] = 1'b0 ^~ inbuffer_data[174];
assign xnor9[175] = 1'b0 ^~ inbuffer_data[175];
assign xnor9[176] = 1'b0 ^~ inbuffer_data[176];
assign xnor9[177] = 1'b0 ^~ inbuffer_data[177];
assign xnor9[178] = 1'b0 ^~ inbuffer_data[178];
assign xnor9[179] = 1'b0 ^~ inbuffer_data[179];
assign xnor9[180] = 1'b1 ^~ inbuffer_data[180];
assign xnor9[181] = 1'b1 ^~ inbuffer_data[181];
assign xnor9[182] = 1'b1 ^~ inbuffer_data[182];
assign xnor9[183] = 1'b1 ^~ inbuffer_data[183];
assign xnor9[184] = 1'b1 ^~ inbuffer_data[184];
assign xnor9[185] = 1'b1 ^~ inbuffer_data[185];
assign xnor9[186] = 1'b1 ^~ inbuffer_data[186];
assign xnor9[187] = 1'b0 ^~ inbuffer_data[187];
assign xnor9[188] = 1'b1 ^~ inbuffer_data[188];
assign xnor9[189] = 1'b0 ^~ inbuffer_data[189];
assign xnor9[190] = 1'b0 ^~ inbuffer_data[190];
assign xnor9[191] = 1'b0 ^~ inbuffer_data[191];
assign xnor9[192] = 1'b0 ^~ inbuffer_data[192];
assign xnor9[193] = 1'b0 ^~ inbuffer_data[193];
assign xnor9[194] = 1'b1 ^~ inbuffer_data[194];
assign xnor9[195] = 1'b0 ^~ inbuffer_data[195];
assign xnor9[196] = 1'b1 ^~ inbuffer_data[196];
assign xnor9[197] = 1'b1 ^~ inbuffer_data[197];
assign xnor9[198] = 1'b1 ^~ inbuffer_data[198];
assign xnor9[199] = 1'b1 ^~ inbuffer_data[199];
assign xnor9[200] = 1'b0 ^~ inbuffer_data[200];
assign xnor9[201] = 1'b0 ^~ inbuffer_data[201];
assign xnor9[202] = 1'b0 ^~ inbuffer_data[202];
assign xnor9[203] = 1'b0 ^~ inbuffer_data[203];
assign xnor9[204] = 1'b0 ^~ inbuffer_data[204];
assign xnor9[205] = 1'b1 ^~ inbuffer_data[205];
assign xnor9[206] = 1'b0 ^~ inbuffer_data[206];
assign xnor9[207] = 1'b1 ^~ inbuffer_data[207];
assign xnor9[208] = 1'b1 ^~ inbuffer_data[208];
assign xnor9[209] = 1'b1 ^~ inbuffer_data[209];
assign xnor9[210] = 1'b1 ^~ inbuffer_data[210];
assign xnor9[211] = 1'b1 ^~ inbuffer_data[211];
assign xnor9[212] = 1'b1 ^~ inbuffer_data[212];
assign xnor9[213] = 1'b1 ^~ inbuffer_data[213];
assign xnor9[214] = 1'b1 ^~ inbuffer_data[214];
assign xnor9[215] = 1'b0 ^~ inbuffer_data[215];
assign xnor9[216] = 1'b1 ^~ inbuffer_data[216];
assign xnor9[217] = 1'b1 ^~ inbuffer_data[217];
assign xnor9[218] = 1'b0 ^~ inbuffer_data[218];
assign xnor9[219] = 1'b0 ^~ inbuffer_data[219];
assign xnor9[220] = 1'b0 ^~ inbuffer_data[220];
assign xnor9[221] = 1'b0 ^~ inbuffer_data[221];
assign xnor9[222] = 1'b0 ^~ inbuffer_data[222];
assign xnor9[223] = 1'b0 ^~ inbuffer_data[223];
assign xnor9[224] = 1'b0 ^~ inbuffer_data[224];
assign xnor9[225] = 1'b1 ^~ inbuffer_data[225];
assign xnor9[226] = 1'b1 ^~ inbuffer_data[226];
assign xnor9[227] = 1'b1 ^~ inbuffer_data[227];
assign xnor9[228] = 1'b0 ^~ inbuffer_data[228];
assign xnor9[229] = 1'b0 ^~ inbuffer_data[229];
assign xnor9[230] = 1'b0 ^~ inbuffer_data[230];
assign xnor9[231] = 1'b0 ^~ inbuffer_data[231];
assign xnor9[232] = 1'b1 ^~ inbuffer_data[232];
assign xnor9[233] = 1'b0 ^~ inbuffer_data[233];
assign xnor9[234] = 1'b0 ^~ inbuffer_data[234];
assign xnor9[235] = 1'b0 ^~ inbuffer_data[235];
assign xnor9[236] = 1'b1 ^~ inbuffer_data[236];
assign xnor9[237] = 1'b1 ^~ inbuffer_data[237];
assign xnor9[238] = 1'b1 ^~ inbuffer_data[238];
assign xnor9[239] = 1'b1 ^~ inbuffer_data[239];
assign xnor9[240] = 1'b1 ^~ inbuffer_data[240];
assign xnor9[241] = 1'b0 ^~ inbuffer_data[241];
assign xnor9[242] = 1'b0 ^~ inbuffer_data[242];
assign xnor9[243] = 1'b1 ^~ inbuffer_data[243];
assign xnor9[244] = 1'b0 ^~ inbuffer_data[244];
assign xnor9[245] = 1'b1 ^~ inbuffer_data[245];
assign xnor9[246] = 1'b0 ^~ inbuffer_data[246];
assign xnor9[247] = 1'b0 ^~ inbuffer_data[247];
assign xnor9[248] = 1'b0 ^~ inbuffer_data[248];
assign xnor9[249] = 1'b0 ^~ inbuffer_data[249];
assign xnor9[250] = 1'b0 ^~ inbuffer_data[250];
assign xnor9[251] = 1'b1 ^~ inbuffer_data[251];
assign xnor9[252] = 1'b1 ^~ inbuffer_data[252];
assign xnor9[253] = 1'b0 ^~ inbuffer_data[253];
assign xnor9[254] = 1'b1 ^~ inbuffer_data[254];
assign xnor9[255] = 1'b0 ^~ inbuffer_data[255];
assign xnor9[256] = 1'b0 ^~ inbuffer_data[256];
assign xnor9[257] = 1'b0 ^~ inbuffer_data[257];
assign xnor9[258] = 1'b1 ^~ inbuffer_data[258];
assign xnor9[259] = 1'b1 ^~ inbuffer_data[259];
assign xnor9[260] = 1'b0 ^~ inbuffer_data[260];
assign xnor9[261] = 1'b0 ^~ inbuffer_data[261];
assign xnor9[262] = 1'b1 ^~ inbuffer_data[262];
assign xnor9[263] = 1'b1 ^~ inbuffer_data[263];
assign xnor9[264] = 1'b1 ^~ inbuffer_data[264];
assign xnor9[265] = 1'b1 ^~ inbuffer_data[265];
assign xnor9[266] = 1'b1 ^~ inbuffer_data[266];
assign xnor9[267] = 1'b1 ^~ inbuffer_data[267];
assign xnor9[268] = 1'b1 ^~ inbuffer_data[268];
assign xnor9[269] = 1'b1 ^~ inbuffer_data[269];
assign xnor9[270] = 1'b1 ^~ inbuffer_data[270];
assign xnor9[271] = 1'b0 ^~ inbuffer_data[271];
assign xnor9[272] = 1'b1 ^~ inbuffer_data[272];
assign xnor9[273] = 1'b0 ^~ inbuffer_data[273];
assign xnor9[274] = 1'b0 ^~ inbuffer_data[274];
assign xnor9[275] = 1'b0 ^~ inbuffer_data[275];
assign xnor9[276] = 1'b0 ^~ inbuffer_data[276];
assign xnor9[277] = 1'b0 ^~ inbuffer_data[277];
assign xnor9[278] = 1'b1 ^~ inbuffer_data[278];
assign xnor9[279] = 1'b1 ^~ inbuffer_data[279];
assign xnor9[280] = 1'b1 ^~ inbuffer_data[280];
assign xnor9[281] = 1'b0 ^~ inbuffer_data[281];
assign xnor9[282] = 1'b1 ^~ inbuffer_data[282];
assign xnor9[283] = 1'b0 ^~ inbuffer_data[283];
assign xnor9[284] = 1'b0 ^~ inbuffer_data[284];
assign xnor9[285] = 1'b1 ^~ inbuffer_data[285];
assign xnor9[286] = 1'b1 ^~ inbuffer_data[286];
assign xnor9[287] = 1'b1 ^~ inbuffer_data[287];
assign xnor9[288] = 1'b1 ^~ inbuffer_data[288];
assign xnor9[289] = 1'b1 ^~ inbuffer_data[289];
assign xnor9[290] = 1'b1 ^~ inbuffer_data[290];
assign xnor9[291] = 1'b1 ^~ inbuffer_data[291];
assign xnor9[292] = 1'b1 ^~ inbuffer_data[292];
assign xnor9[293] = 1'b0 ^~ inbuffer_data[293];
assign xnor9[294] = 1'b0 ^~ inbuffer_data[294];
assign xnor9[295] = 1'b0 ^~ inbuffer_data[295];
assign xnor9[296] = 1'b0 ^~ inbuffer_data[296];
assign xnor9[297] = 1'b1 ^~ inbuffer_data[297];
assign xnor9[298] = 1'b0 ^~ inbuffer_data[298];
assign xnor9[299] = 1'b1 ^~ inbuffer_data[299];
assign xnor9[300] = 1'b1 ^~ inbuffer_data[300];
assign xnor9[301] = 1'b0 ^~ inbuffer_data[301];
assign xnor9[302] = 1'b1 ^~ inbuffer_data[302];
assign xnor9[303] = 1'b0 ^~ inbuffer_data[303];
assign xnor9[304] = 1'b0 ^~ inbuffer_data[304];
assign xnor9[305] = 1'b0 ^~ inbuffer_data[305];
assign xnor9[306] = 1'b0 ^~ inbuffer_data[306];
assign xnor9[307] = 1'b1 ^~ inbuffer_data[307];
assign xnor9[308] = 1'b1 ^~ inbuffer_data[308];
assign xnor9[309] = 1'b0 ^~ inbuffer_data[309];
assign xnor9[310] = 1'b1 ^~ inbuffer_data[310];
assign xnor9[311] = 1'b0 ^~ inbuffer_data[311];
assign xnor9[312] = 1'b0 ^~ inbuffer_data[312];
assign xnor9[313] = 1'b1 ^~ inbuffer_data[313];
assign xnor9[314] = 1'b1 ^~ inbuffer_data[314];
assign xnor9[315] = 1'b1 ^~ inbuffer_data[315];
assign xnor9[316] = 1'b1 ^~ inbuffer_data[316];
assign xnor9[317] = 1'b1 ^~ inbuffer_data[317];
assign xnor9[318] = 1'b1 ^~ inbuffer_data[318];
assign xnor9[319] = 1'b1 ^~ inbuffer_data[319];
assign xnor9[320] = 1'b1 ^~ inbuffer_data[320];
assign xnor9[321] = 1'b0 ^~ inbuffer_data[321];
assign xnor9[322] = 1'b0 ^~ inbuffer_data[322];
assign xnor9[323] = 1'b1 ^~ inbuffer_data[323];
assign xnor9[324] = 1'b1 ^~ inbuffer_data[324];
assign xnor9[325] = 1'b1 ^~ inbuffer_data[325];
assign xnor9[326] = 1'b1 ^~ inbuffer_data[326];
assign xnor9[327] = 1'b1 ^~ inbuffer_data[327];
assign xnor9[328] = 1'b1 ^~ inbuffer_data[328];
assign xnor9[329] = 1'b1 ^~ inbuffer_data[329];
assign xnor9[330] = 1'b1 ^~ inbuffer_data[330];
assign xnor9[331] = 1'b0 ^~ inbuffer_data[331];
assign xnor9[332] = 1'b0 ^~ inbuffer_data[332];
assign xnor9[333] = 1'b0 ^~ inbuffer_data[333];
assign xnor9[334] = 1'b1 ^~ inbuffer_data[334];
assign xnor9[335] = 1'b0 ^~ inbuffer_data[335];
assign xnor9[336] = 1'b0 ^~ inbuffer_data[336];
assign xnor9[337] = 1'b1 ^~ inbuffer_data[337];
assign xnor9[338] = 1'b0 ^~ inbuffer_data[338];
assign xnor9[339] = 1'b0 ^~ inbuffer_data[339];
assign xnor9[340] = 1'b1 ^~ inbuffer_data[340];
assign xnor9[341] = 1'b1 ^~ inbuffer_data[341];
assign xnor9[342] = 1'b1 ^~ inbuffer_data[342];
assign xnor9[343] = 1'b1 ^~ inbuffer_data[343];
assign xnor9[344] = 1'b1 ^~ inbuffer_data[344];
assign xnor9[345] = 1'b1 ^~ inbuffer_data[345];
assign xnor9[346] = 1'b1 ^~ inbuffer_data[346];
assign xnor9[347] = 1'b1 ^~ inbuffer_data[347];
assign xnor9[348] = 1'b0 ^~ inbuffer_data[348];
assign xnor9[349] = 1'b1 ^~ inbuffer_data[349];
assign xnor9[350] = 1'b1 ^~ inbuffer_data[350];
assign xnor9[351] = 1'b1 ^~ inbuffer_data[351];
assign xnor9[352] = 1'b1 ^~ inbuffer_data[352];
assign xnor9[353] = 1'b1 ^~ inbuffer_data[353];
assign xnor9[354] = 1'b1 ^~ inbuffer_data[354];
assign xnor9[355] = 1'b1 ^~ inbuffer_data[355];
assign xnor9[356] = 1'b1 ^~ inbuffer_data[356];
assign xnor9[357] = 1'b1 ^~ inbuffer_data[357];
assign xnor9[358] = 1'b1 ^~ inbuffer_data[358];
assign xnor9[359] = 1'b0 ^~ inbuffer_data[359];
assign xnor9[360] = 1'b1 ^~ inbuffer_data[360];
assign xnor9[361] = 1'b0 ^~ inbuffer_data[361];
assign xnor9[362] = 1'b0 ^~ inbuffer_data[362];
assign xnor9[363] = 1'b0 ^~ inbuffer_data[363];
assign xnor9[364] = 1'b1 ^~ inbuffer_data[364];
assign xnor9[365] = 1'b1 ^~ inbuffer_data[365];
assign xnor9[366] = 1'b1 ^~ inbuffer_data[366];
assign xnor9[367] = 1'b0 ^~ inbuffer_data[367];
assign xnor9[368] = 1'b1 ^~ inbuffer_data[368];
assign xnor9[369] = 1'b1 ^~ inbuffer_data[369];
assign xnor9[370] = 1'b1 ^~ inbuffer_data[370];
assign xnor9[371] = 1'b1 ^~ inbuffer_data[371];
assign xnor9[372] = 1'b1 ^~ inbuffer_data[372];
assign xnor9[373] = 1'b0 ^~ inbuffer_data[373];
assign xnor9[374] = 1'b1 ^~ inbuffer_data[374];
assign xnor9[375] = 1'b1 ^~ inbuffer_data[375];
assign xnor9[376] = 1'b0 ^~ inbuffer_data[376];
assign xnor9[377] = 1'b1 ^~ inbuffer_data[377];
assign xnor9[378] = 1'b1 ^~ inbuffer_data[378];
assign xnor9[379] = 1'b1 ^~ inbuffer_data[379];
assign xnor9[380] = 1'b1 ^~ inbuffer_data[380];
assign xnor9[381] = 1'b1 ^~ inbuffer_data[381];
assign xnor9[382] = 1'b1 ^~ inbuffer_data[382];
assign xnor9[383] = 1'b1 ^~ inbuffer_data[383];
assign xnor9[384] = 1'b1 ^~ inbuffer_data[384];
assign xnor9[385] = 1'b1 ^~ inbuffer_data[385];
assign xnor9[386] = 1'b1 ^~ inbuffer_data[386];
assign xnor9[387] = 1'b0 ^~ inbuffer_data[387];
assign xnor9[388] = 1'b0 ^~ inbuffer_data[388];
assign xnor9[389] = 1'b1 ^~ inbuffer_data[389];
assign xnor9[390] = 1'b0 ^~ inbuffer_data[390];
assign xnor9[391] = 1'b0 ^~ inbuffer_data[391];
assign xnor9[392] = 1'b1 ^~ inbuffer_data[392];
assign xnor9[393] = 1'b1 ^~ inbuffer_data[393];
assign xnor9[394] = 1'b1 ^~ inbuffer_data[394];
assign xnor9[395] = 1'b1 ^~ inbuffer_data[395];
assign xnor9[396] = 1'b1 ^~ inbuffer_data[396];
assign xnor9[397] = 1'b1 ^~ inbuffer_data[397];
assign xnor9[398] = 1'b1 ^~ inbuffer_data[398];
assign xnor9[399] = 1'b1 ^~ inbuffer_data[399];
assign xnor9[400] = 1'b1 ^~ inbuffer_data[400];
assign xnor9[401] = 1'b0 ^~ inbuffer_data[401];
assign xnor9[402] = 1'b0 ^~ inbuffer_data[402];
assign xnor9[403] = 1'b1 ^~ inbuffer_data[403];
assign xnor9[404] = 1'b0 ^~ inbuffer_data[404];
assign xnor9[405] = 1'b1 ^~ inbuffer_data[405];
assign xnor9[406] = 1'b1 ^~ inbuffer_data[406];
assign xnor9[407] = 1'b1 ^~ inbuffer_data[407];
assign xnor9[408] = 1'b1 ^~ inbuffer_data[408];
assign xnor9[409] = 1'b1 ^~ inbuffer_data[409];
assign xnor9[410] = 1'b1 ^~ inbuffer_data[410];
assign xnor9[411] = 1'b1 ^~ inbuffer_data[411];
assign xnor9[412] = 1'b1 ^~ inbuffer_data[412];
assign xnor9[413] = 1'b1 ^~ inbuffer_data[413];
assign xnor9[414] = 1'b1 ^~ inbuffer_data[414];
assign xnor9[415] = 1'b0 ^~ inbuffer_data[415];
assign xnor9[416] = 1'b0 ^~ inbuffer_data[416];
assign xnor9[417] = 1'b1 ^~ inbuffer_data[417];
assign xnor9[418] = 1'b1 ^~ inbuffer_data[418];
assign xnor9[419] = 1'b1 ^~ inbuffer_data[419];
assign xnor9[420] = 1'b1 ^~ inbuffer_data[420];
assign xnor9[421] = 1'b1 ^~ inbuffer_data[421];
assign xnor9[422] = 1'b0 ^~ inbuffer_data[422];
assign xnor9[423] = 1'b1 ^~ inbuffer_data[423];
assign xnor9[424] = 1'b1 ^~ inbuffer_data[424];
assign xnor9[425] = 1'b1 ^~ inbuffer_data[425];
assign xnor9[426] = 1'b1 ^~ inbuffer_data[426];
assign xnor9[427] = 1'b0 ^~ inbuffer_data[427];
assign xnor9[428] = 1'b1 ^~ inbuffer_data[428];
assign xnor9[429] = 1'b1 ^~ inbuffer_data[429];
assign xnor9[430] = 1'b0 ^~ inbuffer_data[430];
assign xnor9[431] = 1'b0 ^~ inbuffer_data[431];
assign xnor9[432] = 1'b0 ^~ inbuffer_data[432];
assign xnor9[433] = 1'b0 ^~ inbuffer_data[433];
assign xnor9[434] = 1'b0 ^~ inbuffer_data[434];
assign xnor9[435] = 1'b1 ^~ inbuffer_data[435];
assign xnor9[436] = 1'b1 ^~ inbuffer_data[436];
assign xnor9[437] = 1'b1 ^~ inbuffer_data[437];
assign xnor9[438] = 1'b1 ^~ inbuffer_data[438];
assign xnor9[439] = 1'b0 ^~ inbuffer_data[439];
assign xnor9[440] = 1'b1 ^~ inbuffer_data[440];
assign xnor9[441] = 1'b1 ^~ inbuffer_data[441];
assign xnor9[442] = 1'b0 ^~ inbuffer_data[442];
assign xnor9[443] = 1'b0 ^~ inbuffer_data[443];
assign xnor9[444] = 1'b0 ^~ inbuffer_data[444];
assign xnor9[445] = 1'b0 ^~ inbuffer_data[445];
assign xnor9[446] = 1'b0 ^~ inbuffer_data[446];
assign xnor9[447] = 1'b1 ^~ inbuffer_data[447];
assign xnor9[448] = 1'b0 ^~ inbuffer_data[448];
assign xnor9[449] = 1'b0 ^~ inbuffer_data[449];
assign xnor9[450] = 1'b0 ^~ inbuffer_data[450];
assign xnor9[451] = 1'b0 ^~ inbuffer_data[451];
assign xnor9[452] = 1'b1 ^~ inbuffer_data[452];
assign xnor9[453] = 1'b1 ^~ inbuffer_data[453];
assign xnor9[454] = 1'b1 ^~ inbuffer_data[454];
assign xnor9[455] = 1'b0 ^~ inbuffer_data[455];
assign xnor9[456] = 1'b1 ^~ inbuffer_data[456];
assign xnor9[457] = 1'b1 ^~ inbuffer_data[457];
assign xnor9[458] = 1'b1 ^~ inbuffer_data[458];
assign xnor9[459] = 1'b1 ^~ inbuffer_data[459];
assign xnor9[460] = 1'b1 ^~ inbuffer_data[460];
assign xnor9[461] = 1'b0 ^~ inbuffer_data[461];
assign xnor9[462] = 1'b0 ^~ inbuffer_data[462];
assign xnor9[463] = 1'b1 ^~ inbuffer_data[463];
assign xnor9[464] = 1'b1 ^~ inbuffer_data[464];
assign xnor9[465] = 1'b1 ^~ inbuffer_data[465];
assign xnor9[466] = 1'b0 ^~ inbuffer_data[466];
assign xnor9[467] = 1'b0 ^~ inbuffer_data[467];
assign xnor9[468] = 1'b1 ^~ inbuffer_data[468];
assign xnor9[469] = 1'b0 ^~ inbuffer_data[469];
assign xnor9[470] = 1'b0 ^~ inbuffer_data[470];
assign xnor9[471] = 1'b0 ^~ inbuffer_data[471];
assign xnor9[472] = 1'b0 ^~ inbuffer_data[472];
assign xnor9[473] = 1'b1 ^~ inbuffer_data[473];
assign xnor9[474] = 1'b0 ^~ inbuffer_data[474];
assign xnor9[475] = 1'b1 ^~ inbuffer_data[475];
assign xnor9[476] = 1'b1 ^~ inbuffer_data[476];
assign xnor9[477] = 1'b1 ^~ inbuffer_data[477];
assign xnor9[478] = 1'b0 ^~ inbuffer_data[478];
assign xnor9[479] = 1'b1 ^~ inbuffer_data[479];
assign xnor9[480] = 1'b0 ^~ inbuffer_data[480];
assign xnor9[481] = 1'b0 ^~ inbuffer_data[481];
assign xnor9[482] = 1'b0 ^~ inbuffer_data[482];
assign xnor9[483] = 1'b1 ^~ inbuffer_data[483];
assign xnor9[484] = 1'b1 ^~ inbuffer_data[484];
assign xnor9[485] = 1'b1 ^~ inbuffer_data[485];
assign xnor9[486] = 1'b1 ^~ inbuffer_data[486];
assign xnor9[487] = 1'b1 ^~ inbuffer_data[487];
assign xnor9[488] = 1'b1 ^~ inbuffer_data[488];
assign xnor9[489] = 1'b0 ^~ inbuffer_data[489];
assign xnor9[490] = 1'b1 ^~ inbuffer_data[490];
assign xnor9[491] = 1'b1 ^~ inbuffer_data[491];
assign xnor9[492] = 1'b0 ^~ inbuffer_data[492];
assign xnor9[493] = 1'b1 ^~ inbuffer_data[493];
assign xnor9[494] = 1'b0 ^~ inbuffer_data[494];
assign xnor9[495] = 1'b0 ^~ inbuffer_data[495];
assign xnor9[496] = 1'b0 ^~ inbuffer_data[496];
assign xnor9[497] = 1'b0 ^~ inbuffer_data[497];
assign xnor9[498] = 1'b0 ^~ inbuffer_data[498];
assign xnor9[499] = 1'b0 ^~ inbuffer_data[499];
assign xnor9[500] = 1'b0 ^~ inbuffer_data[500];
assign xnor9[501] = 1'b1 ^~ inbuffer_data[501];
assign xnor9[502] = 1'b0 ^~ inbuffer_data[502];
assign xnor9[503] = 1'b0 ^~ inbuffer_data[503];
assign xnor9[504] = 1'b0 ^~ inbuffer_data[504];
assign xnor9[505] = 1'b0 ^~ inbuffer_data[505];
assign xnor9[506] = 1'b1 ^~ inbuffer_data[506];
assign xnor9[507] = 1'b0 ^~ inbuffer_data[507];
assign xnor9[508] = 1'b0 ^~ inbuffer_data[508];
assign xnor9[509] = 1'b0 ^~ inbuffer_data[509];
assign xnor9[510] = 1'b1 ^~ inbuffer_data[510];
assign xnor9[511] = 1'b0 ^~ inbuffer_data[511];
assign xnor9[512] = 1'b1 ^~ inbuffer_data[512];
assign xnor9[513] = 1'b0 ^~ inbuffer_data[513];
assign xnor9[514] = 1'b0 ^~ inbuffer_data[514];
assign xnor9[515] = 1'b1 ^~ inbuffer_data[515];
assign xnor9[516] = 1'b0 ^~ inbuffer_data[516];
assign xnor9[517] = 1'b0 ^~ inbuffer_data[517];
assign xnor9[518] = 1'b1 ^~ inbuffer_data[518];
assign xnor9[519] = 1'b0 ^~ inbuffer_data[519];
assign xnor9[520] = 1'b1 ^~ inbuffer_data[520];
assign xnor9[521] = 1'b1 ^~ inbuffer_data[521];
assign xnor9[522] = 1'b0 ^~ inbuffer_data[522];
assign xnor9[523] = 1'b1 ^~ inbuffer_data[523];
assign xnor9[524] = 1'b0 ^~ inbuffer_data[524];
assign xnor9[525] = 1'b0 ^~ inbuffer_data[525];
assign xnor9[526] = 1'b0 ^~ inbuffer_data[526];
assign xnor9[527] = 1'b0 ^~ inbuffer_data[527];
assign xnor9[528] = 1'b0 ^~ inbuffer_data[528];
assign xnor9[529] = 1'b0 ^~ inbuffer_data[529];
assign xnor9[530] = 1'b1 ^~ inbuffer_data[530];
assign xnor9[531] = 1'b1 ^~ inbuffer_data[531];
assign xnor9[532] = 1'b1 ^~ inbuffer_data[532];
assign xnor9[533] = 1'b0 ^~ inbuffer_data[533];
assign xnor9[534] = 1'b0 ^~ inbuffer_data[534];
assign xnor9[535] = 1'b1 ^~ inbuffer_data[535];
assign xnor9[536] = 1'b0 ^~ inbuffer_data[536];
assign xnor9[537] = 1'b0 ^~ inbuffer_data[537];
assign xnor9[538] = 1'b0 ^~ inbuffer_data[538];
assign xnor9[539] = 1'b0 ^~ inbuffer_data[539];
assign xnor9[540] = 1'b0 ^~ inbuffer_data[540];
assign xnor9[541] = 1'b0 ^~ inbuffer_data[541];
assign xnor9[542] = 1'b0 ^~ inbuffer_data[542];
assign xnor9[543] = 1'b0 ^~ inbuffer_data[543];
assign xnor9[544] = 1'b0 ^~ inbuffer_data[544];
assign xnor9[545] = 1'b0 ^~ inbuffer_data[545];
assign xnor9[546] = 1'b1 ^~ inbuffer_data[546];
assign xnor9[547] = 1'b0 ^~ inbuffer_data[547];
assign xnor9[548] = 1'b0 ^~ inbuffer_data[548];
assign xnor9[549] = 1'b0 ^~ inbuffer_data[549];
assign xnor9[550] = 1'b0 ^~ inbuffer_data[550];
assign xnor9[551] = 1'b1 ^~ inbuffer_data[551];
assign xnor9[552] = 1'b1 ^~ inbuffer_data[552];
assign xnor9[553] = 1'b0 ^~ inbuffer_data[553];
assign xnor9[554] = 1'b0 ^~ inbuffer_data[554];
assign xnor9[555] = 1'b0 ^~ inbuffer_data[555];
assign xnor9[556] = 1'b1 ^~ inbuffer_data[556];
assign xnor9[557] = 1'b0 ^~ inbuffer_data[557];
assign xnor9[558] = 1'b1 ^~ inbuffer_data[558];
assign xnor9[559] = 1'b0 ^~ inbuffer_data[559];
assign xnor9[560] = 1'b1 ^~ inbuffer_data[560];
assign xnor9[561] = 1'b1 ^~ inbuffer_data[561];
assign xnor9[562] = 1'b0 ^~ inbuffer_data[562];
assign xnor9[563] = 1'b0 ^~ inbuffer_data[563];
assign xnor9[564] = 1'b1 ^~ inbuffer_data[564];
assign xnor9[565] = 1'b0 ^~ inbuffer_data[565];
assign xnor9[566] = 1'b0 ^~ inbuffer_data[566];
assign xnor9[567] = 1'b0 ^~ inbuffer_data[567];
assign xnor9[568] = 1'b0 ^~ inbuffer_data[568];
assign xnor9[569] = 1'b0 ^~ inbuffer_data[569];
assign xnor9[570] = 1'b0 ^~ inbuffer_data[570];
assign xnor9[571] = 1'b0 ^~ inbuffer_data[571];
assign xnor9[572] = 1'b0 ^~ inbuffer_data[572];
assign xnor9[573] = 1'b0 ^~ inbuffer_data[573];
assign xnor9[574] = 1'b0 ^~ inbuffer_data[574];
assign xnor9[575] = 1'b0 ^~ inbuffer_data[575];
assign xnor9[576] = 1'b0 ^~ inbuffer_data[576];
assign xnor9[577] = 1'b1 ^~ inbuffer_data[577];
assign xnor9[578] = 1'b0 ^~ inbuffer_data[578];
assign xnor9[579] = 1'b1 ^~ inbuffer_data[579];
assign xnor9[580] = 1'b1 ^~ inbuffer_data[580];
assign xnor9[581] = 1'b0 ^~ inbuffer_data[581];
assign xnor9[582] = 1'b0 ^~ inbuffer_data[582];
assign xnor9[583] = 1'b1 ^~ inbuffer_data[583];
assign xnor9[584] = 1'b0 ^~ inbuffer_data[584];
assign xnor9[585] = 1'b1 ^~ inbuffer_data[585];
assign xnor9[586] = 1'b1 ^~ inbuffer_data[586];
assign xnor9[587] = 1'b1 ^~ inbuffer_data[587];
assign xnor9[588] = 1'b1 ^~ inbuffer_data[588];
assign xnor9[589] = 1'b0 ^~ inbuffer_data[589];
assign xnor9[590] = 1'b1 ^~ inbuffer_data[590];
assign xnor9[591] = 1'b0 ^~ inbuffer_data[591];
assign xnor9[592] = 1'b1 ^~ inbuffer_data[592];
assign xnor9[593] = 1'b0 ^~ inbuffer_data[593];
assign xnor9[594] = 1'b1 ^~ inbuffer_data[594];
assign xnor9[595] = 1'b0 ^~ inbuffer_data[595];
assign xnor9[596] = 1'b0 ^~ inbuffer_data[596];
assign xnor9[597] = 1'b0 ^~ inbuffer_data[597];
assign xnor9[598] = 1'b0 ^~ inbuffer_data[598];
assign xnor9[599] = 1'b0 ^~ inbuffer_data[599];
assign xnor9[600] = 1'b0 ^~ inbuffer_data[600];
assign xnor9[601] = 1'b0 ^~ inbuffer_data[601];
assign xnor9[602] = 1'b0 ^~ inbuffer_data[602];
assign xnor9[603] = 1'b0 ^~ inbuffer_data[603];
assign xnor9[604] = 1'b0 ^~ inbuffer_data[604];
assign xnor9[605] = 1'b0 ^~ inbuffer_data[605];
assign xnor9[606] = 1'b0 ^~ inbuffer_data[606];
assign xnor9[607] = 1'b0 ^~ inbuffer_data[607];
assign xnor9[608] = 1'b1 ^~ inbuffer_data[608];
assign xnor9[609] = 1'b1 ^~ inbuffer_data[609];
assign xnor9[610] = 1'b0 ^~ inbuffer_data[610];
assign xnor9[611] = 1'b0 ^~ inbuffer_data[611];
assign xnor9[612] = 1'b1 ^~ inbuffer_data[612];
assign xnor9[613] = 1'b1 ^~ inbuffer_data[613];
assign xnor9[614] = 1'b0 ^~ inbuffer_data[614];
assign xnor9[615] = 1'b1 ^~ inbuffer_data[615];
assign xnor9[616] = 1'b0 ^~ inbuffer_data[616];
assign xnor9[617] = 1'b0 ^~ inbuffer_data[617];
assign xnor9[618] = 1'b1 ^~ inbuffer_data[618];
assign xnor9[619] = 1'b1 ^~ inbuffer_data[619];
assign xnor9[620] = 1'b0 ^~ inbuffer_data[620];
assign xnor9[621] = 1'b0 ^~ inbuffer_data[621];
assign xnor9[622] = 1'b0 ^~ inbuffer_data[622];
assign xnor9[623] = 1'b0 ^~ inbuffer_data[623];
assign xnor9[624] = 1'b0 ^~ inbuffer_data[624];
assign xnor9[625] = 1'b1 ^~ inbuffer_data[625];
assign xnor9[626] = 1'b0 ^~ inbuffer_data[626];
assign xnor9[627] = 1'b1 ^~ inbuffer_data[627];
assign xnor9[628] = 1'b0 ^~ inbuffer_data[628];
assign xnor9[629] = 1'b0 ^~ inbuffer_data[629];
assign xnor9[630] = 1'b0 ^~ inbuffer_data[630];
assign xnor9[631] = 1'b0 ^~ inbuffer_data[631];
assign xnor9[632] = 1'b0 ^~ inbuffer_data[632];
assign xnor9[633] = 1'b0 ^~ inbuffer_data[633];
assign xnor9[634] = 1'b1 ^~ inbuffer_data[634];
assign xnor9[635] = 1'b0 ^~ inbuffer_data[635];
assign xnor9[636] = 1'b0 ^~ inbuffer_data[636];
assign xnor9[637] = 1'b0 ^~ inbuffer_data[637];
assign xnor9[638] = 1'b1 ^~ inbuffer_data[638];
assign xnor9[639] = 1'b1 ^~ inbuffer_data[639];
assign xnor9[640] = 1'b0 ^~ inbuffer_data[640];
assign xnor9[641] = 1'b1 ^~ inbuffer_data[641];
assign xnor9[642] = 1'b1 ^~ inbuffer_data[642];
assign xnor9[643] = 1'b0 ^~ inbuffer_data[643];
assign xnor9[644] = 1'b0 ^~ inbuffer_data[644];
assign xnor9[645] = 1'b1 ^~ inbuffer_data[645];
assign xnor9[646] = 1'b0 ^~ inbuffer_data[646];
assign xnor9[647] = 1'b0 ^~ inbuffer_data[647];
assign xnor9[648] = 1'b0 ^~ inbuffer_data[648];
assign xnor9[649] = 1'b0 ^~ inbuffer_data[649];
assign xnor9[650] = 1'b0 ^~ inbuffer_data[650];
assign xnor9[651] = 1'b0 ^~ inbuffer_data[651];
assign xnor9[652] = 1'b1 ^~ inbuffer_data[652];
assign xnor9[653] = 1'b0 ^~ inbuffer_data[653];
assign xnor9[654] = 1'b0 ^~ inbuffer_data[654];
assign xnor9[655] = 1'b0 ^~ inbuffer_data[655];
assign xnor9[656] = 1'b1 ^~ inbuffer_data[656];
assign xnor9[657] = 1'b1 ^~ inbuffer_data[657];
assign xnor9[658] = 1'b0 ^~ inbuffer_data[658];
assign xnor9[659] = 1'b0 ^~ inbuffer_data[659];
assign xnor9[660] = 1'b0 ^~ inbuffer_data[660];
assign xnor9[661] = 1'b0 ^~ inbuffer_data[661];
assign xnor9[662] = 1'b0 ^~ inbuffer_data[662];
assign xnor9[663] = 1'b0 ^~ inbuffer_data[663];
assign xnor9[664] = 1'b1 ^~ inbuffer_data[664];
assign xnor9[665] = 1'b1 ^~ inbuffer_data[665];
assign xnor9[666] = 1'b1 ^~ inbuffer_data[666];
assign xnor9[667] = 1'b0 ^~ inbuffer_data[667];
assign xnor9[668] = 1'b0 ^~ inbuffer_data[668];
assign xnor9[669] = 1'b0 ^~ inbuffer_data[669];
assign xnor9[670] = 1'b0 ^~ inbuffer_data[670];
assign xnor9[671] = 1'b0 ^~ inbuffer_data[671];
assign xnor9[672] = 1'b0 ^~ inbuffer_data[672];
assign xnor9[673] = 1'b0 ^~ inbuffer_data[673];
assign xnor9[674] = 1'b1 ^~ inbuffer_data[674];
assign xnor9[675] = 1'b1 ^~ inbuffer_data[675];
assign xnor9[676] = 1'b0 ^~ inbuffer_data[676];
assign xnor9[677] = 1'b0 ^~ inbuffer_data[677];
assign xnor9[678] = 1'b1 ^~ inbuffer_data[678];
assign xnor9[679] = 1'b1 ^~ inbuffer_data[679];
assign xnor9[680] = 1'b1 ^~ inbuffer_data[680];
assign xnor9[681] = 1'b0 ^~ inbuffer_data[681];
assign xnor9[682] = 1'b1 ^~ inbuffer_data[682];
assign xnor9[683] = 1'b0 ^~ inbuffer_data[683];
assign xnor9[684] = 1'b0 ^~ inbuffer_data[684];
assign xnor9[685] = 1'b0 ^~ inbuffer_data[685];
assign xnor9[686] = 1'b1 ^~ inbuffer_data[686];
assign xnor9[687] = 1'b0 ^~ inbuffer_data[687];
assign xnor9[688] = 1'b1 ^~ inbuffer_data[688];
assign xnor9[689] = 1'b1 ^~ inbuffer_data[689];
assign xnor9[690] = 1'b1 ^~ inbuffer_data[690];
assign xnor9[691] = 1'b1 ^~ inbuffer_data[691];
assign xnor9[692] = 1'b1 ^~ inbuffer_data[692];
assign xnor9[693] = 1'b1 ^~ inbuffer_data[693];
assign xnor9[694] = 1'b1 ^~ inbuffer_data[694];
assign xnor9[695] = 1'b1 ^~ inbuffer_data[695];
assign xnor9[696] = 1'b0 ^~ inbuffer_data[696];
assign xnor9[697] = 1'b0 ^~ inbuffer_data[697];
assign xnor9[698] = 1'b1 ^~ inbuffer_data[698];
assign xnor9[699] = 1'b0 ^~ inbuffer_data[699];
assign xnor9[700] = 1'b0 ^~ inbuffer_data[700];
assign xnor9[701] = 1'b1 ^~ inbuffer_data[701];
assign xnor9[702] = 1'b0 ^~ inbuffer_data[702];
assign xnor9[703] = 1'b1 ^~ inbuffer_data[703];
assign xnor9[704] = 1'b0 ^~ inbuffer_data[704];
assign xnor9[705] = 1'b1 ^~ inbuffer_data[705];
assign xnor9[706] = 1'b0 ^~ inbuffer_data[706];
assign xnor9[707] = 1'b1 ^~ inbuffer_data[707];
assign xnor9[708] = 1'b1 ^~ inbuffer_data[708];
assign xnor9[709] = 1'b1 ^~ inbuffer_data[709];
assign xnor9[710] = 1'b1 ^~ inbuffer_data[710];
assign xnor9[711] = 1'b1 ^~ inbuffer_data[711];
assign xnor9[712] = 1'b1 ^~ inbuffer_data[712];
assign xnor9[713] = 1'b1 ^~ inbuffer_data[713];
assign xnor9[714] = 1'b1 ^~ inbuffer_data[714];
assign xnor9[715] = 1'b1 ^~ inbuffer_data[715];
assign xnor9[716] = 1'b1 ^~ inbuffer_data[716];
assign xnor9[717] = 1'b1 ^~ inbuffer_data[717];
assign xnor9[718] = 1'b1 ^~ inbuffer_data[718];
assign xnor9[719] = 1'b1 ^~ inbuffer_data[719];
assign xnor9[720] = 1'b1 ^~ inbuffer_data[720];
assign xnor9[721] = 1'b1 ^~ inbuffer_data[721];
assign xnor9[722] = 1'b1 ^~ inbuffer_data[722];
assign xnor9[723] = 1'b0 ^~ inbuffer_data[723];
assign xnor9[724] = 1'b0 ^~ inbuffer_data[724];
assign xnor9[725] = 1'b0 ^~ inbuffer_data[725];
assign xnor9[726] = 1'b0 ^~ inbuffer_data[726];
assign xnor9[727] = 1'b1 ^~ inbuffer_data[727];
assign xnor9[728] = 1'b1 ^~ inbuffer_data[728];
assign xnor9[729] = 1'b1 ^~ inbuffer_data[729];
assign xnor9[730] = 1'b1 ^~ inbuffer_data[730];
assign xnor9[731] = 1'b1 ^~ inbuffer_data[731];
assign xnor9[732] = 1'b1 ^~ inbuffer_data[732];
assign xnor9[733] = 1'b0 ^~ inbuffer_data[733];
assign xnor9[734] = 1'b0 ^~ inbuffer_data[734];
assign xnor9[735] = 1'b1 ^~ inbuffer_data[735];
assign xnor9[736] = 1'b1 ^~ inbuffer_data[736];
assign xnor9[737] = 1'b1 ^~ inbuffer_data[737];
assign xnor9[738] = 1'b1 ^~ inbuffer_data[738];
assign xnor9[739] = 1'b1 ^~ inbuffer_data[739];
assign xnor9[740] = 1'b1 ^~ inbuffer_data[740];
assign xnor9[741] = 1'b1 ^~ inbuffer_data[741];
assign xnor9[742] = 1'b1 ^~ inbuffer_data[742];
assign xnor9[743] = 1'b1 ^~ inbuffer_data[743];
assign xnor9[744] = 1'b1 ^~ inbuffer_data[744];
assign xnor9[745] = 1'b1 ^~ inbuffer_data[745];
assign xnor9[746] = 1'b1 ^~ inbuffer_data[746];
assign xnor9[747] = 1'b1 ^~ inbuffer_data[747];
assign xnor9[748] = 1'b1 ^~ inbuffer_data[748];
assign xnor9[749] = 1'b1 ^~ inbuffer_data[749];
assign xnor9[750] = 1'b1 ^~ inbuffer_data[750];
assign xnor9[751] = 1'b0 ^~ inbuffer_data[751];
assign xnor9[752] = 1'b1 ^~ inbuffer_data[752];
assign xnor9[753] = 1'b1 ^~ inbuffer_data[753];
assign xnor9[754] = 1'b1 ^~ inbuffer_data[754];
assign xnor9[755] = 1'b0 ^~ inbuffer_data[755];
assign xnor9[756] = 1'b0 ^~ inbuffer_data[756];
assign xnor9[757] = 1'b1 ^~ inbuffer_data[757];
assign xnor9[758] = 1'b0 ^~ inbuffer_data[758];
assign xnor9[759] = 1'b0 ^~ inbuffer_data[759];
assign xnor9[760] = 1'b0 ^~ inbuffer_data[760];
assign xnor9[761] = 1'b0 ^~ inbuffer_data[761];
assign xnor9[762] = 1'b0 ^~ inbuffer_data[762];
assign xnor9[763] = 1'b0 ^~ inbuffer_data[763];
assign xnor9[764] = 1'b1 ^~ inbuffer_data[764];
assign xnor9[765] = 1'b1 ^~ inbuffer_data[765];
assign xnor9[766] = 1'b0 ^~ inbuffer_data[766];
assign xnor9[767] = 1'b0 ^~ inbuffer_data[767];
assign xnor9[768] = 1'b1 ^~ inbuffer_data[768];
assign xnor9[769] = 1'b0 ^~ inbuffer_data[769];
assign xnor9[770] = 1'b1 ^~ inbuffer_data[770];
assign xnor9[771] = 1'b1 ^~ inbuffer_data[771];
assign xnor9[772] = 1'b0 ^~ inbuffer_data[772];
assign xnor9[773] = 1'b0 ^~ inbuffer_data[773];
assign xnor9[774] = 1'b0 ^~ inbuffer_data[774];
assign xnor9[775] = 1'b0 ^~ inbuffer_data[775];
assign xnor9[776] = 1'b1 ^~ inbuffer_data[776];
assign xnor9[777] = 1'b0 ^~ inbuffer_data[777];
assign xnor9[778] = 1'b1 ^~ inbuffer_data[778];
assign xnor9[779] = 1'b0 ^~ inbuffer_data[779];
assign xnor9[780] = 1'b0 ^~ inbuffer_data[780];
assign xnor9[781] = 1'b1 ^~ inbuffer_data[781];
assign xnor9[782] = 1'b0 ^~ inbuffer_data[782];
assign xnor9[783] = 1'b0 ^~ inbuffer_data[783];

endmodule