module layer_0_conv #(
    parameter INPUT_DIM = 28,   //28x28
    parameter OUTPUT_DIM = 10,
    parameter KERNEL_DIM = 3,
    parameter INPUT_CHANNELS = 1,
    parameter OUTPUT_CHANNELS = 2,
    parameter DATATYPE_SIZE = 1
) (
    input clk,
    input reset,

    input i_we,
    input [DATATYPE_SIZE-1:0] i_data [INPUT_CHANNELS-1:0],

    output [DATATYPE_SIZE-1:0] o_data [OUTPUT_CHANNELS-1:0],
    output o_we
);

localparam TEMP_SIZE = INPUT_CHANNELS * OUTPUT_CHANNELS * (KERNAL_DIM ** 2);

reg window [INPUT_CHANNELS-1:0][KERNAL_DIM**2-1:0];
reg temp [TEMP_SIZE-1:0];

ibuf_conv #(
                        .img_width(INPUT_DIM),
                        .kernel_dim(KERNEL_DIM),
                    ) ibuf (
                        .clk(clk),
                        .i_we(i_we),
                        .i_data(i_data[0]),
                        .o_data(window[0]),
                    );

# ibuf_conv #(
#     .img_width(INPUT_DIM),
#     .kernel_dim(KERNEL_DIM),
# ) ibuf (
#     .clk(clk),
#     .i_we(i_we),
#     .i_data(i_data[%INPUT_C%]),
#     .o_data(window[%INPUT_C%]),
# );

assign temp[0] = ~window[0][0];
assign temp[1] = ~window[0][1];
assign temp[2] = ~window[0][2];
assign temp[3] = ~window[0][3];
assign temp[4] = window[0][4];
assign temp[5] = ~window[0][5];
assign temp[6] = window[0][6];
assign temp[7] = ~window[0][7];
assign temp[8] = window[0][8];
assign temp[9] = window[0][9];
assign temp[10] = window[0][10];
assign temp[11] = ~window[0][11];
assign temp[12] = window[0][12];
assign temp[13] = window[0][13];
assign temp[14] = window[0][14];
assign temp[15] = ~window[0][15];
assign temp[32] = ~window[0][0];
assign temp[33] = ~window[0][1];
assign temp[34] = ~window[0][2];
assign temp[35] = ~window[0][3];
assign temp[36] = ~window[0][4];
assign temp[37] = ~window[0][5];
assign temp[38] = window[0][6];
assign temp[39] = ~window[0][7];
assign temp[40] = window[0][8];
assign temp[41] = window[0][9];
assign temp[42] = window[0][10];
assign temp[43] = ~window[0][11];
assign temp[44] = window[0][12];
assign temp[45] = window[0][13];
assign temp[46] = window[0][14];
assign temp[47] = ~window[0][15];
assign temp[64] = ~window[0][0];
assign temp[65] = window[0][1];
assign temp[66] = ~window[0][2];
assign temp[67] = ~window[0][3];
assign temp[68] = ~window[0][4];
assign temp[69] = ~window[0][5];
assign temp[70] = ~window[0][6];
assign temp[71] = ~window[0][7];
assign temp[72] = ~window[0][8];
assign temp[73] = ~window[0][9];
assign temp[74] = ~window[0][10];
assign temp[75] = window[0][11];
assign temp[76] = window[0][12];
assign temp[77] = window[0][13];
assign temp[78] = window[0][14];
assign temp[79] = window[0][15];
assign temp[96] = window[0][0];
assign temp[97] = window[0][1];
assign temp[98] = ~window[0][2];
assign temp[99] = ~window[0][3];
assign temp[100] = window[0][4];
assign temp[101] = ~window[0][5];
assign temp[102] = ~window[0][6];
assign temp[103] = ~window[0][7];
assign temp[104] = window[0][8];
assign temp[105] = ~window[0][9];
assign temp[106] = ~window[0][10];
assign temp[107] = ~window[0][11];
assign temp[108] = window[0][12];
assign temp[109] = ~window[0][13];
assign temp[110] = ~window[0][14];
assign temp[111] = ~window[0][15];
assign temp[128] = window[0][0];
assign temp[129] = window[0][1];
assign temp[130] = ~window[0][2];
assign temp[131] = ~window[0][3];
assign temp[132] = window[0][4];
assign temp[133] = ~window[0][5];
assign temp[134] = ~window[0][6];
assign temp[135] = window[0][7];
assign temp[136] = window[0][8];
assign temp[137] = window[0][9];
assign temp[138] = window[0][10];
assign temp[139] = window[0][11];
assign temp[140] = window[0][12];
assign temp[141] = window[0][13];
assign temp[142] = window[0][14];
assign temp[143] = ~window[0][15];
assign temp[160] = ~window[0][0];
assign temp[161] = window[0][1];
assign temp[162] = window[0][2];
assign temp[163] = window[0][3];
assign temp[164] = ~window[0][4];
assign temp[165] = ~window[0][5];
assign temp[166] = window[0][6];
assign temp[167] = window[0][7];
assign temp[168] = ~window[0][8];
assign temp[169] = ~window[0][9];
assign temp[170] = ~window[0][10];
assign temp[171] = ~window[0][11];
assign temp[172] = ~window[0][12];
assign temp[173] = ~window[0][13];
assign temp[174] = window[0][14];
assign temp[175] = window[0][15];
assign temp[192] = ~window[0][0];
assign temp[193] = window[0][1];
assign temp[194] = window[0][2];
assign temp[195] = window[0][3];
assign temp[196] = ~window[0][4];
assign temp[197] = ~window[0][5];
assign temp[198] = ~window[0][6];
assign temp[199] = ~window[0][7];
assign temp[200] = ~window[0][8];
assign temp[201] = ~window[0][9];
assign temp[202] = ~window[0][10];
assign temp[203] = ~window[0][11];
assign temp[204] = ~window[0][12];
assign temp[205] = ~window[0][13];
assign temp[206] = ~window[0][14];
assign temp[207] = ~window[0][15];
assign temp[224] = ~window[0][0];
assign temp[225] = ~window[0][1];
assign temp[226] = ~window[0][2];
assign temp[227] = ~window[0][3];
assign temp[228] = ~window[0][4];
assign temp[229] = ~window[0][5];
assign temp[230] = ~window[0][6];
assign temp[231] = ~window[0][7];
assign temp[232] = ~window[0][8];
assign temp[233] = ~window[0][9];
assign temp[234] = ~window[0][10];
assign temp[235] = ~window[0][11];
assign temp[236] = window[0][12];
assign temp[237] = window[0][13];
assign temp[238] = window[0][14];
assign temp[239] = window[0][15];
assign temp[256] = ~window[0][0];
assign temp[257] = ~window[0][1];
assign temp[258] = window[0][2];
assign temp[259] = window[0][3];
assign temp[260] = window[0][4];
assign temp[261] = window[0][5];
assign temp[262] = window[0][6];
assign temp[263] = window[0][7];
assign temp[264] = ~window[0][8];
assign temp[265] = window[0][9];
assign temp[266] = window[0][10];
assign temp[267] = window[0][11];
assign temp[268] = ~window[0][12];
assign temp[269] = ~window[0][13];
assign temp[270] = ~window[0][14];
assign temp[271] = window[0][15];
assign temp[288] = ~window[0][0];
assign temp[289] = ~window[0][1];
assign temp[290] = ~window[0][2];
assign temp[291] = window[0][3];
assign temp[292] = ~window[0][4];
assign temp[293] = ~window[0][5];
assign temp[294] = ~window[0][6];
assign temp[295] = window[0][7];
assign temp[296] = ~window[0][8];
assign temp[297] = ~window[0][9];
assign temp[298] = ~window[0][10];
assign temp[299] = window[0][11];
assign temp[300] = window[0][12];
assign temp[301] = window[0][13];
assign temp[302] = window[0][14];
assign temp[303] = window[0][15];
assign temp[320] = window[0][0];
assign temp[321] = window[0][1];
assign temp[322] = window[0][2];
assign temp[323] = window[0][3];
assign temp[324] = window[0][4];
assign temp[325] = window[0][5];
assign temp[326] = ~window[0][6];
assign temp[327] = ~window[0][7];
assign temp[328] = window[0][8];
assign temp[329] = window[0][9];
assign temp[330] = ~window[0][10];
assign temp[331] = window[0][11];
assign temp[332] = window[0][12];
assign temp[333] = window[0][13];
assign temp[334] = window[0][14];
assign temp[335] = ~window[0][15];
assign temp[352] = ~window[0][0];
assign temp[353] = ~window[0][1];
assign temp[354] = window[0][2];
assign temp[355] = window[0][3];
assign temp[356] = ~window[0][4];
assign temp[357] = ~window[0][5];
assign temp[358] = ~window[0][6];
assign temp[359] = ~window[0][7];
assign temp[360] = ~window[0][8];
assign temp[361] = ~window[0][9];
assign temp[362] = ~window[0][10];
assign temp[363] = ~window[0][11];
assign temp[364] = window[0][12];
assign temp[365] = ~window[0][13];
assign temp[366] = window[0][14];
assign temp[367] = ~window[0][15];
assign temp[384] = ~window[0][0];
assign temp[385] = window[0][1];
assign temp[386] = ~window[0][2];
assign temp[387] = ~window[0][3];
assign temp[388] = window[0][4];
assign temp[389] = ~window[0][5];
assign temp[390] = ~window[0][6];
assign temp[391] = ~window[0][7];
assign temp[392] = ~window[0][8];
assign temp[393] = ~window[0][9];
assign temp[394] = ~window[0][10];
assign temp[395] = window[0][11];
assign temp[396] = ~window[0][12];
assign temp[397] = ~window[0][13];
assign temp[398] = ~window[0][14];
assign temp[399] = window[0][15];
assign temp[416] = ~window[0][0];
assign temp[417] = ~window[0][1];
assign temp[418] = ~window[0][2];
assign temp[419] = ~window[0][3];
assign temp[420] = ~window[0][4];
assign temp[421] = window[0][5];
assign temp[422] = window[0][6];
assign temp[423] = window[0][7];
assign temp[424] = window[0][8];
assign temp[425] = window[0][9];
assign temp[426] = window[0][10];
assign temp[427] = ~window[0][11];
assign temp[428] = ~window[0][12];
assign temp[429] = ~window[0][13];
assign temp[430] = window[0][14];
assign temp[431] = window[0][15];
assign temp[448] = window[0][0];
assign temp[449] = window[0][1];
assign temp[450] = ~window[0][2];
assign temp[451] = window[0][3];
assign temp[452] = window[0][4];
assign temp[453] = window[0][5];
assign temp[454] = window[0][6];
assign temp[455] = window[0][7];
assign temp[456] = window[0][8];
assign temp[457] = window[0][9];
assign temp[458] = window[0][10];
assign temp[459] = ~window[0][11];
assign temp[460] = ~window[0][12];
assign temp[461] = ~window[0][13];
assign temp[462] = ~window[0][14];
assign temp[463] = ~window[0][15];
assign temp[480] = ~window[0][0];
assign temp[481] = window[0][1];
assign temp[482] = window[0][2];
assign temp[483] = window[0][3];
assign temp[484] = window[0][4];
assign temp[485] = window[0][5];
assign temp[486] = ~window[0][6];
assign temp[487] = ~window[0][7];
assign temp[488] = window[0][8];
assign temp[489] = ~window[0][9];
assign temp[490] = ~window[0][10];
assign temp[491] = ~window[0][11];
assign temp[492] = window[0][12];
assign temp[493] = window[0][13];
assign temp[494] = ~window[0][14];
assign temp[495] = ~window[0][15];
assign temp[512] = window[0][0];
assign temp[513] = window[0][1];
assign temp[514] = ~window[0][2];
assign temp[515] = window[0][3];
assign temp[516] = window[0][4];
assign temp[517] = ~window[0][5];
assign temp[518] = window[0][6];
assign temp[519] = window[0][7];
assign temp[520] = window[0][8];
assign temp[521] = ~window[0][9];
assign temp[522] = window[0][10];
assign temp[523] = window[0][11];
assign temp[524] = window[0][12];
assign temp[525] = ~window[0][13];
assign temp[526] = window[0][14];
assign temp[527] = window[0][15];
assign temp[544] = ~window[0][0];
assign temp[545] = ~window[0][1];
assign temp[546] = window[0][2];
assign temp[547] = window[0][3];
assign temp[548] = ~window[0][4];
assign temp[549] = ~window[0][5];
assign temp[550] = window[0][6];
assign temp[551] = window[0][7];
assign temp[552] = window[0][8];
assign temp[553] = window[0][9];
assign temp[554] = ~window[0][10];
assign temp[555] = window[0][11];
assign temp[556] = ~window[0][12];
assign temp[557] = window[0][13];
assign temp[558] = window[0][14];
assign temp[559] = window[0][15];
assign temp[576] = ~window[0][0];
assign temp[577] = ~window[0][1];
assign temp[578] = ~window[0][2];
assign temp[579] = window[0][3];
assign temp[580] = ~window[0][4];
assign temp[581] = ~window[0][5];
assign temp[582] = ~window[0][6];
assign temp[583] = ~window[0][7];
assign temp[584] = window[0][8];
assign temp[585] = window[0][9];
assign temp[586] = ~window[0][10];
assign temp[587] = ~window[0][11];
assign temp[588] = window[0][12];
assign temp[589] = window[0][13];
assign temp[590] = window[0][14];
assign temp[591] = window[0][15];
assign temp[608] = ~window[0][0];
assign temp[609] = window[0][1];
assign temp[610] = window[0][2];
assign temp[611] = window[0][3];
assign temp[612] = window[0][4];
assign temp[613] = window[0][5];
assign temp[614] = ~window[0][6];
assign temp[615] = ~window[0][7];
assign temp[616] = window[0][8];
assign temp[617] = ~window[0][9];
assign temp[618] = ~window[0][10];
assign temp[619] = ~window[0][11];
assign temp[620] = ~window[0][12];
assign temp[621] = window[0][13];
assign temp[622] = ~window[0][14];
assign temp[623] = ~window[0][15];
assign temp[640] = ~window[0][0];
assign temp[641] = ~window[0][1];
assign temp[642] = ~window[0][2];
assign temp[643] = ~window[0][3];
assign temp[644] = ~window[0][4];
assign temp[645] = ~window[0][5];
assign temp[646] = ~window[0][6];
assign temp[647] = ~window[0][7];
assign temp[648] = ~window[0][8];
assign temp[649] = ~window[0][9];
assign temp[650] = window[0][10];
assign temp[651] = window[0][11];
assign temp[652] = ~window[0][12];
assign temp[653] = window[0][13];
assign temp[654] = window[0][14];
assign temp[655] = window[0][15];
assign temp[672] = ~window[0][0];
assign temp[673] = window[0][1];
assign temp[674] = ~window[0][2];
assign temp[675] = window[0][3];
assign temp[676] = window[0][4];
assign temp[677] = window[0][5];
assign temp[678] = ~window[0][6];
assign temp[679] = window[0][7];
assign temp[680] = window[0][8];
assign temp[681] = window[0][9];
assign temp[682] = ~window[0][10];
assign temp[683] = window[0][11];
assign temp[684] = window[0][12];
assign temp[685] = window[0][13];
assign temp[686] = ~window[0][14];
assign temp[687] = ~window[0][15];
assign temp[704] = ~window[0][0];
assign temp[705] = ~window[0][1];
assign temp[706] = ~window[0][2];
assign temp[707] = ~window[0][3];
assign temp[708] = ~window[0][4];
assign temp[709] = window[0][5];
assign temp[710] = ~window[0][6];
assign temp[711] = ~window[0][7];
assign temp[712] = window[0][8];
assign temp[713] = window[0][9];
assign temp[714] = window[0][10];
assign temp[715] = window[0][11];
assign temp[716] = window[0][12];
assign temp[717] = window[0][13];
assign temp[718] = window[0][14];
assign temp[719] = window[0][15];
assign temp[736] = ~window[0][0];
assign temp[737] = ~window[0][1];
assign temp[738] = ~window[0][2];
assign temp[739] = ~window[0][3];
assign temp[740] = window[0][4];
assign temp[741] = window[0][5];
assign temp[742] = window[0][6];
assign temp[743] = ~window[0][7];
assign temp[744] = window[0][8];
assign temp[745] = window[0][9];
assign temp[746] = window[0][10];
assign temp[747] = ~window[0][11];
assign temp[748] = window[0][12];
assign temp[749] = ~window[0][13];
assign temp[750] = ~window[0][14];
assign temp[751] = window[0][15];
assign temp[768] = window[0][0];
assign temp[769] = ~window[0][1];
assign temp[770] = ~window[0][2];
assign temp[771] = window[0][3];
assign temp[772] = ~window[0][4];
assign temp[773] = ~window[0][5];
assign temp[774] = ~window[0][6];
assign temp[775] = ~window[0][7];
assign temp[776] = window[0][8];
assign temp[777] = window[0][9];
assign temp[778] = ~window[0][10];
assign temp[779] = ~window[0][11];
assign temp[780] = window[0][12];
assign temp[781] = window[0][13];
assign temp[782] = window[0][14];
assign temp[783] = ~window[0][15];
assign temp[800] = window[0][0];
assign temp[801] = ~window[0][1];
assign temp[802] = window[0][2];
assign temp[803] = ~window[0][3];
assign temp[804] = window[0][4];
assign temp[805] = window[0][5];
assign temp[806] = ~window[0][6];
assign temp[807] = window[0][7];
assign temp[808] = ~window[0][8];
assign temp[809] = ~window[0][9];
assign temp[810] = ~window[0][10];
assign temp[811] = window[0][11];
assign temp[812] = ~window[0][12];
assign temp[813] = ~window[0][13];
assign temp[814] = ~window[0][14];
assign temp[815] = window[0][15];
assign temp[832] = window[0][0];
assign temp[833] = window[0][1];
assign temp[834] = window[0][2];
assign temp[835] = window[0][3];
assign temp[836] = ~window[0][4];
assign temp[837] = ~window[0][5];
assign temp[838] = window[0][6];
assign temp[839] = window[0][7];
assign temp[840] = ~window[0][8];
assign temp[841] = ~window[0][9];
assign temp[842] = ~window[0][10];
assign temp[843] = ~window[0][11];
assign temp[844] = ~window[0][12];
assign temp[845] = ~window[0][13];
assign temp[846] = ~window[0][14];
assign temp[847] = ~window[0][15];
assign temp[864] = ~window[0][0];
assign temp[865] = ~window[0][1];
assign temp[866] = ~window[0][2];
assign temp[867] = ~window[0][3];
assign temp[868] = ~window[0][4];
assign temp[869] = ~window[0][5];
assign temp[870] = ~window[0][6];
assign temp[871] = ~window[0][7];
assign temp[872] = ~window[0][8];
assign temp[873] = ~window[0][9];
assign temp[874] = ~window[0][10];
assign temp[875] = ~window[0][11];
assign temp[876] = ~window[0][12];
assign temp[877] = ~window[0][13];
assign temp[878] = ~window[0][14];
assign temp[879] = window[0][15];
assign temp[896] = window[0][0];
assign temp[897] = window[0][1];
assign temp[898] = window[0][2];
assign temp[899] = ~window[0][3];
assign temp[900] = window[0][4];
assign temp[901] = window[0][5];
assign temp[902] = ~window[0][6];
assign temp[903] = ~window[0][7];
assign temp[904] = window[0][8];
assign temp[905] = window[0][9];
assign temp[906] = ~window[0][10];
assign temp[907] = ~window[0][11];
assign temp[908] = window[0][12];
assign temp[909] = ~window[0][13];
assign temp[910] = ~window[0][14];
assign temp[911] = ~window[0][15];
assign temp[928] = ~window[0][0];
assign temp[929] = ~window[0][1];
assign temp[930] = window[0][2];
assign temp[931] = window[0][3];
assign temp[932] = window[0][4];
assign temp[933] = window[0][5];
assign temp[934] = window[0][6];
assign temp[935] = window[0][7];
assign temp[936] = ~window[0][8];
assign temp[937] = window[0][9];
assign temp[938] = ~window[0][10];
assign temp[939] = ~window[0][11];
assign temp[940] = ~window[0][12];
assign temp[941] = window[0][13];
assign temp[942] = window[0][14];
assign temp[943] = ~window[0][15];
assign temp[960] = window[0][0];
assign temp[961] = ~window[0][1];
assign temp[962] = ~window[0][2];
assign temp[963] = ~window[0][3];
assign temp[964] = ~window[0][4];
assign temp[965] = window[0][5];
assign temp[966] = ~window[0][6];
assign temp[967] = ~window[0][7];
assign temp[968] = window[0][8];
assign temp[969] = window[0][9];
assign temp[970] = window[0][10];
assign temp[971] = ~window[0][11];
assign temp[972] = window[0][12];
assign temp[973] = window[0][13];
assign temp[974] = ~window[0][14];
assign temp[975] = ~window[0][15];
assign temp[992] = ~window[0][0];
assign temp[993] = ~window[0][1];
assign temp[994] = window[0][2];
assign temp[995] = ~window[0][3];
assign temp[996] = ~window[0][4];
assign temp[997] = window[0][5];
assign temp[998] = window[0][6];
assign temp[999] = ~window[0][7];
assign temp[1000] = window[0][8];
assign temp[1001] = window[0][9];
assign temp[1002] = window[0][10];
assign temp[1003] = window[0][11];
assign temp[1004] = window[0][12];
assign temp[1005] = window[0][13];
assign temp[1006] = window[0][14];
assign temp[1007] = window[0][15];


always @(*) begin
    for (int i = 0; i < OUTPUT_CHANNELS; i++) begin
        for (int j = 0; j < INPUT_CHANNELS; j++) begin
            for (int k = 0; k < KERNEL_DIM ** 2; k++) begin
            o[i] += temp[i * OUTPUT_CHANNELS + j * INPUT_CHANNELS + k];
            end
        end
    end
end
endmodule